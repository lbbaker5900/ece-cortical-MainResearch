
            begin
              gen[0][0].run()  ;
            end
            begin
              drv[0][0].run()  ;
            end
            begin
              dma2mem[0][0].run()  ;
            end

            begin
              gen[0][1].run()  ;
            end
            begin
              drv[0][1].run()  ;
            end
            begin
              dma2mem[0][1].run()  ;
            end

            begin
              gen[0][2].run()  ;
            end
            begin
              drv[0][2].run()  ;
            end
            begin
              dma2mem[0][2].run()  ;
            end

            begin
              gen[0][3].run()  ;
            end
            begin
              drv[0][3].run()  ;
            end
            begin
              dma2mem[0][3].run()  ;
            end

            begin
              gen[0][4].run()  ;
            end
            begin
              drv[0][4].run()  ;
            end
            begin
              dma2mem[0][4].run()  ;
            end

            begin
              gen[0][5].run()  ;
            end
            begin
              drv[0][5].run()  ;
            end
            begin
              dma2mem[0][5].run()  ;
            end

            begin
              gen[0][6].run()  ;
            end
            begin
              drv[0][6].run()  ;
            end
            begin
              dma2mem[0][6].run()  ;
            end

            begin
              gen[0][7].run()  ;
            end
            begin
              drv[0][7].run()  ;
            end
            begin
              dma2mem[0][7].run()  ;
            end

            begin
              gen[0][8].run()  ;
            end
            begin
              drv[0][8].run()  ;
            end
            begin
              dma2mem[0][8].run()  ;
            end

            begin
              gen[0][9].run()  ;
            end
            begin
              drv[0][9].run()  ;
            end
            begin
              dma2mem[0][9].run()  ;
            end

            begin
              gen[0][10].run()  ;
            end
            begin
              drv[0][10].run()  ;
            end
            begin
              dma2mem[0][10].run()  ;
            end

            begin
              gen[0][11].run()  ;
            end
            begin
              drv[0][11].run()  ;
            end
            begin
              dma2mem[0][11].run()  ;
            end

            begin
              gen[0][12].run()  ;
            end
            begin
              drv[0][12].run()  ;
            end
            begin
              dma2mem[0][12].run()  ;
            end

            begin
              gen[0][13].run()  ;
            end
            begin
              drv[0][13].run()  ;
            end
            begin
              dma2mem[0][13].run()  ;
            end

            begin
              gen[0][14].run()  ;
            end
            begin
              drv[0][14].run()  ;
            end
            begin
              dma2mem[0][14].run()  ;
            end

            begin
              gen[0][15].run()  ;
            end
            begin
              drv[0][15].run()  ;
            end
            begin
              dma2mem[0][15].run()  ;
            end

            begin
              gen[0][16].run()  ;
            end
            begin
              drv[0][16].run()  ;
            end
            begin
              dma2mem[0][16].run()  ;
            end

            begin
              gen[0][17].run()  ;
            end
            begin
              drv[0][17].run()  ;
            end
            begin
              dma2mem[0][17].run()  ;
            end

            begin
              gen[0][18].run()  ;
            end
            begin
              drv[0][18].run()  ;
            end
            begin
              dma2mem[0][18].run()  ;
            end

            begin
              gen[0][19].run()  ;
            end
            begin
              drv[0][19].run()  ;
            end
            begin
              dma2mem[0][19].run()  ;
            end

            begin
              gen[0][20].run()  ;
            end
            begin
              drv[0][20].run()  ;
            end
            begin
              dma2mem[0][20].run()  ;
            end

            begin
              gen[0][21].run()  ;
            end
            begin
              drv[0][21].run()  ;
            end
            begin
              dma2mem[0][21].run()  ;
            end

            begin
              gen[0][22].run()  ;
            end
            begin
              drv[0][22].run()  ;
            end
            begin
              dma2mem[0][22].run()  ;
            end

            begin
              gen[0][23].run()  ;
            end
            begin
              drv[0][23].run()  ;
            end
            begin
              dma2mem[0][23].run()  ;
            end

            begin
              gen[0][24].run()  ;
            end
            begin
              drv[0][24].run()  ;
            end
            begin
              dma2mem[0][24].run()  ;
            end

            begin
              gen[0][25].run()  ;
            end
            begin
              drv[0][25].run()  ;
            end
            begin
              dma2mem[0][25].run()  ;
            end

            begin
              gen[0][26].run()  ;
            end
            begin
              drv[0][26].run()  ;
            end
            begin
              dma2mem[0][26].run()  ;
            end

            begin
              gen[0][27].run()  ;
            end
            begin
              drv[0][27].run()  ;
            end
            begin
              dma2mem[0][27].run()  ;
            end

            begin
              gen[0][28].run()  ;
            end
            begin
              drv[0][28].run()  ;
            end
            begin
              dma2mem[0][28].run()  ;
            end

            begin
              gen[0][29].run()  ;
            end
            begin
              drv[0][29].run()  ;
            end
            begin
              dma2mem[0][29].run()  ;
            end

            begin
              gen[0][30].run()  ;
            end
            begin
              drv[0][30].run()  ;
            end
            begin
              dma2mem[0][30].run()  ;
            end

            begin
              gen[0][31].run()  ;
            end
            begin
              drv[0][31].run()  ;
            end
            begin
              dma2mem[0][31].run()  ;
            end

            begin
              gen[1][0].run()  ;
            end
            begin
              drv[1][0].run()  ;
            end
            begin
              dma2mem[1][0].run()  ;
            end

            begin
              gen[1][1].run()  ;
            end
            begin
              drv[1][1].run()  ;
            end
            begin
              dma2mem[1][1].run()  ;
            end

            begin
              gen[1][2].run()  ;
            end
            begin
              drv[1][2].run()  ;
            end
            begin
              dma2mem[1][2].run()  ;
            end

            begin
              gen[1][3].run()  ;
            end
            begin
              drv[1][3].run()  ;
            end
            begin
              dma2mem[1][3].run()  ;
            end

            begin
              gen[1][4].run()  ;
            end
            begin
              drv[1][4].run()  ;
            end
            begin
              dma2mem[1][4].run()  ;
            end

            begin
              gen[1][5].run()  ;
            end
            begin
              drv[1][5].run()  ;
            end
            begin
              dma2mem[1][5].run()  ;
            end

            begin
              gen[1][6].run()  ;
            end
            begin
              drv[1][6].run()  ;
            end
            begin
              dma2mem[1][6].run()  ;
            end

            begin
              gen[1][7].run()  ;
            end
            begin
              drv[1][7].run()  ;
            end
            begin
              dma2mem[1][7].run()  ;
            end

            begin
              gen[1][8].run()  ;
            end
            begin
              drv[1][8].run()  ;
            end
            begin
              dma2mem[1][8].run()  ;
            end

            begin
              gen[1][9].run()  ;
            end
            begin
              drv[1][9].run()  ;
            end
            begin
              dma2mem[1][9].run()  ;
            end

            begin
              gen[1][10].run()  ;
            end
            begin
              drv[1][10].run()  ;
            end
            begin
              dma2mem[1][10].run()  ;
            end

            begin
              gen[1][11].run()  ;
            end
            begin
              drv[1][11].run()  ;
            end
            begin
              dma2mem[1][11].run()  ;
            end

            begin
              gen[1][12].run()  ;
            end
            begin
              drv[1][12].run()  ;
            end
            begin
              dma2mem[1][12].run()  ;
            end

            begin
              gen[1][13].run()  ;
            end
            begin
              drv[1][13].run()  ;
            end
            begin
              dma2mem[1][13].run()  ;
            end

            begin
              gen[1][14].run()  ;
            end
            begin
              drv[1][14].run()  ;
            end
            begin
              dma2mem[1][14].run()  ;
            end

            begin
              gen[1][15].run()  ;
            end
            begin
              drv[1][15].run()  ;
            end
            begin
              dma2mem[1][15].run()  ;
            end

            begin
              gen[1][16].run()  ;
            end
            begin
              drv[1][16].run()  ;
            end
            begin
              dma2mem[1][16].run()  ;
            end

            begin
              gen[1][17].run()  ;
            end
            begin
              drv[1][17].run()  ;
            end
            begin
              dma2mem[1][17].run()  ;
            end

            begin
              gen[1][18].run()  ;
            end
            begin
              drv[1][18].run()  ;
            end
            begin
              dma2mem[1][18].run()  ;
            end

            begin
              gen[1][19].run()  ;
            end
            begin
              drv[1][19].run()  ;
            end
            begin
              dma2mem[1][19].run()  ;
            end

            begin
              gen[1][20].run()  ;
            end
            begin
              drv[1][20].run()  ;
            end
            begin
              dma2mem[1][20].run()  ;
            end

            begin
              gen[1][21].run()  ;
            end
            begin
              drv[1][21].run()  ;
            end
            begin
              dma2mem[1][21].run()  ;
            end

            begin
              gen[1][22].run()  ;
            end
            begin
              drv[1][22].run()  ;
            end
            begin
              dma2mem[1][22].run()  ;
            end

            begin
              gen[1][23].run()  ;
            end
            begin
              drv[1][23].run()  ;
            end
            begin
              dma2mem[1][23].run()  ;
            end

            begin
              gen[1][24].run()  ;
            end
            begin
              drv[1][24].run()  ;
            end
            begin
              dma2mem[1][24].run()  ;
            end

            begin
              gen[1][25].run()  ;
            end
            begin
              drv[1][25].run()  ;
            end
            begin
              dma2mem[1][25].run()  ;
            end

            begin
              gen[1][26].run()  ;
            end
            begin
              drv[1][26].run()  ;
            end
            begin
              dma2mem[1][26].run()  ;
            end

            begin
              gen[1][27].run()  ;
            end
            begin
              drv[1][27].run()  ;
            end
            begin
              dma2mem[1][27].run()  ;
            end

            begin
              gen[1][28].run()  ;
            end
            begin
              drv[1][28].run()  ;
            end
            begin
              dma2mem[1][28].run()  ;
            end

            begin
              gen[1][29].run()  ;
            end
            begin
              drv[1][29].run()  ;
            end
            begin
              dma2mem[1][29].run()  ;
            end

            begin
              gen[1][30].run()  ;
            end
            begin
              drv[1][30].run()  ;
            end
            begin
              dma2mem[1][30].run()  ;
            end

            begin
              gen[1][31].run()  ;
            end
            begin
              drv[1][31].run()  ;
            end
            begin
              dma2mem[1][31].run()  ;
            end

            begin
              gen[2][0].run()  ;
            end
            begin
              drv[2][0].run()  ;
            end
            begin
              dma2mem[2][0].run()  ;
            end

            begin
              gen[2][1].run()  ;
            end
            begin
              drv[2][1].run()  ;
            end
            begin
              dma2mem[2][1].run()  ;
            end

            begin
              gen[2][2].run()  ;
            end
            begin
              drv[2][2].run()  ;
            end
            begin
              dma2mem[2][2].run()  ;
            end

            begin
              gen[2][3].run()  ;
            end
            begin
              drv[2][3].run()  ;
            end
            begin
              dma2mem[2][3].run()  ;
            end

            begin
              gen[2][4].run()  ;
            end
            begin
              drv[2][4].run()  ;
            end
            begin
              dma2mem[2][4].run()  ;
            end

            begin
              gen[2][5].run()  ;
            end
            begin
              drv[2][5].run()  ;
            end
            begin
              dma2mem[2][5].run()  ;
            end

            begin
              gen[2][6].run()  ;
            end
            begin
              drv[2][6].run()  ;
            end
            begin
              dma2mem[2][6].run()  ;
            end

            begin
              gen[2][7].run()  ;
            end
            begin
              drv[2][7].run()  ;
            end
            begin
              dma2mem[2][7].run()  ;
            end

            begin
              gen[2][8].run()  ;
            end
            begin
              drv[2][8].run()  ;
            end
            begin
              dma2mem[2][8].run()  ;
            end

            begin
              gen[2][9].run()  ;
            end
            begin
              drv[2][9].run()  ;
            end
            begin
              dma2mem[2][9].run()  ;
            end

            begin
              gen[2][10].run()  ;
            end
            begin
              drv[2][10].run()  ;
            end
            begin
              dma2mem[2][10].run()  ;
            end

            begin
              gen[2][11].run()  ;
            end
            begin
              drv[2][11].run()  ;
            end
            begin
              dma2mem[2][11].run()  ;
            end

            begin
              gen[2][12].run()  ;
            end
            begin
              drv[2][12].run()  ;
            end
            begin
              dma2mem[2][12].run()  ;
            end

            begin
              gen[2][13].run()  ;
            end
            begin
              drv[2][13].run()  ;
            end
            begin
              dma2mem[2][13].run()  ;
            end

            begin
              gen[2][14].run()  ;
            end
            begin
              drv[2][14].run()  ;
            end
            begin
              dma2mem[2][14].run()  ;
            end

            begin
              gen[2][15].run()  ;
            end
            begin
              drv[2][15].run()  ;
            end
            begin
              dma2mem[2][15].run()  ;
            end

            begin
              gen[2][16].run()  ;
            end
            begin
              drv[2][16].run()  ;
            end
            begin
              dma2mem[2][16].run()  ;
            end

            begin
              gen[2][17].run()  ;
            end
            begin
              drv[2][17].run()  ;
            end
            begin
              dma2mem[2][17].run()  ;
            end

            begin
              gen[2][18].run()  ;
            end
            begin
              drv[2][18].run()  ;
            end
            begin
              dma2mem[2][18].run()  ;
            end

            begin
              gen[2][19].run()  ;
            end
            begin
              drv[2][19].run()  ;
            end
            begin
              dma2mem[2][19].run()  ;
            end

            begin
              gen[2][20].run()  ;
            end
            begin
              drv[2][20].run()  ;
            end
            begin
              dma2mem[2][20].run()  ;
            end

            begin
              gen[2][21].run()  ;
            end
            begin
              drv[2][21].run()  ;
            end
            begin
              dma2mem[2][21].run()  ;
            end

            begin
              gen[2][22].run()  ;
            end
            begin
              drv[2][22].run()  ;
            end
            begin
              dma2mem[2][22].run()  ;
            end

            begin
              gen[2][23].run()  ;
            end
            begin
              drv[2][23].run()  ;
            end
            begin
              dma2mem[2][23].run()  ;
            end

            begin
              gen[2][24].run()  ;
            end
            begin
              drv[2][24].run()  ;
            end
            begin
              dma2mem[2][24].run()  ;
            end

            begin
              gen[2][25].run()  ;
            end
            begin
              drv[2][25].run()  ;
            end
            begin
              dma2mem[2][25].run()  ;
            end

            begin
              gen[2][26].run()  ;
            end
            begin
              drv[2][26].run()  ;
            end
            begin
              dma2mem[2][26].run()  ;
            end

            begin
              gen[2][27].run()  ;
            end
            begin
              drv[2][27].run()  ;
            end
            begin
              dma2mem[2][27].run()  ;
            end

            begin
              gen[2][28].run()  ;
            end
            begin
              drv[2][28].run()  ;
            end
            begin
              dma2mem[2][28].run()  ;
            end

            begin
              gen[2][29].run()  ;
            end
            begin
              drv[2][29].run()  ;
            end
            begin
              dma2mem[2][29].run()  ;
            end

            begin
              gen[2][30].run()  ;
            end
            begin
              drv[2][30].run()  ;
            end
            begin
              dma2mem[2][30].run()  ;
            end

            begin
              gen[2][31].run()  ;
            end
            begin
              drv[2][31].run()  ;
            end
            begin
              dma2mem[2][31].run()  ;
            end

            begin
              gen[3][0].run()  ;
            end
            begin
              drv[3][0].run()  ;
            end
            begin
              dma2mem[3][0].run()  ;
            end

            begin
              gen[3][1].run()  ;
            end
            begin
              drv[3][1].run()  ;
            end
            begin
              dma2mem[3][1].run()  ;
            end

            begin
              gen[3][2].run()  ;
            end
            begin
              drv[3][2].run()  ;
            end
            begin
              dma2mem[3][2].run()  ;
            end

            begin
              gen[3][3].run()  ;
            end
            begin
              drv[3][3].run()  ;
            end
            begin
              dma2mem[3][3].run()  ;
            end

            begin
              gen[3][4].run()  ;
            end
            begin
              drv[3][4].run()  ;
            end
            begin
              dma2mem[3][4].run()  ;
            end

            begin
              gen[3][5].run()  ;
            end
            begin
              drv[3][5].run()  ;
            end
            begin
              dma2mem[3][5].run()  ;
            end

            begin
              gen[3][6].run()  ;
            end
            begin
              drv[3][6].run()  ;
            end
            begin
              dma2mem[3][6].run()  ;
            end

            begin
              gen[3][7].run()  ;
            end
            begin
              drv[3][7].run()  ;
            end
            begin
              dma2mem[3][7].run()  ;
            end

            begin
              gen[3][8].run()  ;
            end
            begin
              drv[3][8].run()  ;
            end
            begin
              dma2mem[3][8].run()  ;
            end

            begin
              gen[3][9].run()  ;
            end
            begin
              drv[3][9].run()  ;
            end
            begin
              dma2mem[3][9].run()  ;
            end

            begin
              gen[3][10].run()  ;
            end
            begin
              drv[3][10].run()  ;
            end
            begin
              dma2mem[3][10].run()  ;
            end

            begin
              gen[3][11].run()  ;
            end
            begin
              drv[3][11].run()  ;
            end
            begin
              dma2mem[3][11].run()  ;
            end

            begin
              gen[3][12].run()  ;
            end
            begin
              drv[3][12].run()  ;
            end
            begin
              dma2mem[3][12].run()  ;
            end

            begin
              gen[3][13].run()  ;
            end
            begin
              drv[3][13].run()  ;
            end
            begin
              dma2mem[3][13].run()  ;
            end

            begin
              gen[3][14].run()  ;
            end
            begin
              drv[3][14].run()  ;
            end
            begin
              dma2mem[3][14].run()  ;
            end

            begin
              gen[3][15].run()  ;
            end
            begin
              drv[3][15].run()  ;
            end
            begin
              dma2mem[3][15].run()  ;
            end

            begin
              gen[3][16].run()  ;
            end
            begin
              drv[3][16].run()  ;
            end
            begin
              dma2mem[3][16].run()  ;
            end

            begin
              gen[3][17].run()  ;
            end
            begin
              drv[3][17].run()  ;
            end
            begin
              dma2mem[3][17].run()  ;
            end

            begin
              gen[3][18].run()  ;
            end
            begin
              drv[3][18].run()  ;
            end
            begin
              dma2mem[3][18].run()  ;
            end

            begin
              gen[3][19].run()  ;
            end
            begin
              drv[3][19].run()  ;
            end
            begin
              dma2mem[3][19].run()  ;
            end

            begin
              gen[3][20].run()  ;
            end
            begin
              drv[3][20].run()  ;
            end
            begin
              dma2mem[3][20].run()  ;
            end

            begin
              gen[3][21].run()  ;
            end
            begin
              drv[3][21].run()  ;
            end
            begin
              dma2mem[3][21].run()  ;
            end

            begin
              gen[3][22].run()  ;
            end
            begin
              drv[3][22].run()  ;
            end
            begin
              dma2mem[3][22].run()  ;
            end

            begin
              gen[3][23].run()  ;
            end
            begin
              drv[3][23].run()  ;
            end
            begin
              dma2mem[3][23].run()  ;
            end

            begin
              gen[3][24].run()  ;
            end
            begin
              drv[3][24].run()  ;
            end
            begin
              dma2mem[3][24].run()  ;
            end

            begin
              gen[3][25].run()  ;
            end
            begin
              drv[3][25].run()  ;
            end
            begin
              dma2mem[3][25].run()  ;
            end

            begin
              gen[3][26].run()  ;
            end
            begin
              drv[3][26].run()  ;
            end
            begin
              dma2mem[3][26].run()  ;
            end

            begin
              gen[3][27].run()  ;
            end
            begin
              drv[3][27].run()  ;
            end
            begin
              dma2mem[3][27].run()  ;
            end

            begin
              gen[3][28].run()  ;
            end
            begin
              drv[3][28].run()  ;
            end
            begin
              dma2mem[3][28].run()  ;
            end

            begin
              gen[3][29].run()  ;
            end
            begin
              drv[3][29].run()  ;
            end
            begin
              dma2mem[3][29].run()  ;
            end

            begin
              gen[3][30].run()  ;
            end
            begin
              drv[3][30].run()  ;
            end
            begin
              dma2mem[3][30].run()  ;
            end

            begin
              gen[3][31].run()  ;
            end
            begin
              drv[3][31].run()  ;
            end
            begin
              dma2mem[3][31].run()  ;
            end

            begin
              gen[4][0].run()  ;
            end
            begin
              drv[4][0].run()  ;
            end
            begin
              dma2mem[4][0].run()  ;
            end

            begin
              gen[4][1].run()  ;
            end
            begin
              drv[4][1].run()  ;
            end
            begin
              dma2mem[4][1].run()  ;
            end

            begin
              gen[4][2].run()  ;
            end
            begin
              drv[4][2].run()  ;
            end
            begin
              dma2mem[4][2].run()  ;
            end

            begin
              gen[4][3].run()  ;
            end
            begin
              drv[4][3].run()  ;
            end
            begin
              dma2mem[4][3].run()  ;
            end

            begin
              gen[4][4].run()  ;
            end
            begin
              drv[4][4].run()  ;
            end
            begin
              dma2mem[4][4].run()  ;
            end

            begin
              gen[4][5].run()  ;
            end
            begin
              drv[4][5].run()  ;
            end
            begin
              dma2mem[4][5].run()  ;
            end

            begin
              gen[4][6].run()  ;
            end
            begin
              drv[4][6].run()  ;
            end
            begin
              dma2mem[4][6].run()  ;
            end

            begin
              gen[4][7].run()  ;
            end
            begin
              drv[4][7].run()  ;
            end
            begin
              dma2mem[4][7].run()  ;
            end

            begin
              gen[4][8].run()  ;
            end
            begin
              drv[4][8].run()  ;
            end
            begin
              dma2mem[4][8].run()  ;
            end

            begin
              gen[4][9].run()  ;
            end
            begin
              drv[4][9].run()  ;
            end
            begin
              dma2mem[4][9].run()  ;
            end

            begin
              gen[4][10].run()  ;
            end
            begin
              drv[4][10].run()  ;
            end
            begin
              dma2mem[4][10].run()  ;
            end

            begin
              gen[4][11].run()  ;
            end
            begin
              drv[4][11].run()  ;
            end
            begin
              dma2mem[4][11].run()  ;
            end

            begin
              gen[4][12].run()  ;
            end
            begin
              drv[4][12].run()  ;
            end
            begin
              dma2mem[4][12].run()  ;
            end

            begin
              gen[4][13].run()  ;
            end
            begin
              drv[4][13].run()  ;
            end
            begin
              dma2mem[4][13].run()  ;
            end

            begin
              gen[4][14].run()  ;
            end
            begin
              drv[4][14].run()  ;
            end
            begin
              dma2mem[4][14].run()  ;
            end

            begin
              gen[4][15].run()  ;
            end
            begin
              drv[4][15].run()  ;
            end
            begin
              dma2mem[4][15].run()  ;
            end

            begin
              gen[4][16].run()  ;
            end
            begin
              drv[4][16].run()  ;
            end
            begin
              dma2mem[4][16].run()  ;
            end

            begin
              gen[4][17].run()  ;
            end
            begin
              drv[4][17].run()  ;
            end
            begin
              dma2mem[4][17].run()  ;
            end

            begin
              gen[4][18].run()  ;
            end
            begin
              drv[4][18].run()  ;
            end
            begin
              dma2mem[4][18].run()  ;
            end

            begin
              gen[4][19].run()  ;
            end
            begin
              drv[4][19].run()  ;
            end
            begin
              dma2mem[4][19].run()  ;
            end

            begin
              gen[4][20].run()  ;
            end
            begin
              drv[4][20].run()  ;
            end
            begin
              dma2mem[4][20].run()  ;
            end

            begin
              gen[4][21].run()  ;
            end
            begin
              drv[4][21].run()  ;
            end
            begin
              dma2mem[4][21].run()  ;
            end

            begin
              gen[4][22].run()  ;
            end
            begin
              drv[4][22].run()  ;
            end
            begin
              dma2mem[4][22].run()  ;
            end

            begin
              gen[4][23].run()  ;
            end
            begin
              drv[4][23].run()  ;
            end
            begin
              dma2mem[4][23].run()  ;
            end

            begin
              gen[4][24].run()  ;
            end
            begin
              drv[4][24].run()  ;
            end
            begin
              dma2mem[4][24].run()  ;
            end

            begin
              gen[4][25].run()  ;
            end
            begin
              drv[4][25].run()  ;
            end
            begin
              dma2mem[4][25].run()  ;
            end

            begin
              gen[4][26].run()  ;
            end
            begin
              drv[4][26].run()  ;
            end
            begin
              dma2mem[4][26].run()  ;
            end

            begin
              gen[4][27].run()  ;
            end
            begin
              drv[4][27].run()  ;
            end
            begin
              dma2mem[4][27].run()  ;
            end

            begin
              gen[4][28].run()  ;
            end
            begin
              drv[4][28].run()  ;
            end
            begin
              dma2mem[4][28].run()  ;
            end

            begin
              gen[4][29].run()  ;
            end
            begin
              drv[4][29].run()  ;
            end
            begin
              dma2mem[4][29].run()  ;
            end

            begin
              gen[4][30].run()  ;
            end
            begin
              drv[4][30].run()  ;
            end
            begin
              dma2mem[4][30].run()  ;
            end

            begin
              gen[4][31].run()  ;
            end
            begin
              drv[4][31].run()  ;
            end
            begin
              dma2mem[4][31].run()  ;
            end

            begin
              gen[5][0].run()  ;
            end
            begin
              drv[5][0].run()  ;
            end
            begin
              dma2mem[5][0].run()  ;
            end

            begin
              gen[5][1].run()  ;
            end
            begin
              drv[5][1].run()  ;
            end
            begin
              dma2mem[5][1].run()  ;
            end

            begin
              gen[5][2].run()  ;
            end
            begin
              drv[5][2].run()  ;
            end
            begin
              dma2mem[5][2].run()  ;
            end

            begin
              gen[5][3].run()  ;
            end
            begin
              drv[5][3].run()  ;
            end
            begin
              dma2mem[5][3].run()  ;
            end

            begin
              gen[5][4].run()  ;
            end
            begin
              drv[5][4].run()  ;
            end
            begin
              dma2mem[5][4].run()  ;
            end

            begin
              gen[5][5].run()  ;
            end
            begin
              drv[5][5].run()  ;
            end
            begin
              dma2mem[5][5].run()  ;
            end

            begin
              gen[5][6].run()  ;
            end
            begin
              drv[5][6].run()  ;
            end
            begin
              dma2mem[5][6].run()  ;
            end

            begin
              gen[5][7].run()  ;
            end
            begin
              drv[5][7].run()  ;
            end
            begin
              dma2mem[5][7].run()  ;
            end

            begin
              gen[5][8].run()  ;
            end
            begin
              drv[5][8].run()  ;
            end
            begin
              dma2mem[5][8].run()  ;
            end

            begin
              gen[5][9].run()  ;
            end
            begin
              drv[5][9].run()  ;
            end
            begin
              dma2mem[5][9].run()  ;
            end

            begin
              gen[5][10].run()  ;
            end
            begin
              drv[5][10].run()  ;
            end
            begin
              dma2mem[5][10].run()  ;
            end

            begin
              gen[5][11].run()  ;
            end
            begin
              drv[5][11].run()  ;
            end
            begin
              dma2mem[5][11].run()  ;
            end

            begin
              gen[5][12].run()  ;
            end
            begin
              drv[5][12].run()  ;
            end
            begin
              dma2mem[5][12].run()  ;
            end

            begin
              gen[5][13].run()  ;
            end
            begin
              drv[5][13].run()  ;
            end
            begin
              dma2mem[5][13].run()  ;
            end

            begin
              gen[5][14].run()  ;
            end
            begin
              drv[5][14].run()  ;
            end
            begin
              dma2mem[5][14].run()  ;
            end

            begin
              gen[5][15].run()  ;
            end
            begin
              drv[5][15].run()  ;
            end
            begin
              dma2mem[5][15].run()  ;
            end

            begin
              gen[5][16].run()  ;
            end
            begin
              drv[5][16].run()  ;
            end
            begin
              dma2mem[5][16].run()  ;
            end

            begin
              gen[5][17].run()  ;
            end
            begin
              drv[5][17].run()  ;
            end
            begin
              dma2mem[5][17].run()  ;
            end

            begin
              gen[5][18].run()  ;
            end
            begin
              drv[5][18].run()  ;
            end
            begin
              dma2mem[5][18].run()  ;
            end

            begin
              gen[5][19].run()  ;
            end
            begin
              drv[5][19].run()  ;
            end
            begin
              dma2mem[5][19].run()  ;
            end

            begin
              gen[5][20].run()  ;
            end
            begin
              drv[5][20].run()  ;
            end
            begin
              dma2mem[5][20].run()  ;
            end

            begin
              gen[5][21].run()  ;
            end
            begin
              drv[5][21].run()  ;
            end
            begin
              dma2mem[5][21].run()  ;
            end

            begin
              gen[5][22].run()  ;
            end
            begin
              drv[5][22].run()  ;
            end
            begin
              dma2mem[5][22].run()  ;
            end

            begin
              gen[5][23].run()  ;
            end
            begin
              drv[5][23].run()  ;
            end
            begin
              dma2mem[5][23].run()  ;
            end

            begin
              gen[5][24].run()  ;
            end
            begin
              drv[5][24].run()  ;
            end
            begin
              dma2mem[5][24].run()  ;
            end

            begin
              gen[5][25].run()  ;
            end
            begin
              drv[5][25].run()  ;
            end
            begin
              dma2mem[5][25].run()  ;
            end

            begin
              gen[5][26].run()  ;
            end
            begin
              drv[5][26].run()  ;
            end
            begin
              dma2mem[5][26].run()  ;
            end

            begin
              gen[5][27].run()  ;
            end
            begin
              drv[5][27].run()  ;
            end
            begin
              dma2mem[5][27].run()  ;
            end

            begin
              gen[5][28].run()  ;
            end
            begin
              drv[5][28].run()  ;
            end
            begin
              dma2mem[5][28].run()  ;
            end

            begin
              gen[5][29].run()  ;
            end
            begin
              drv[5][29].run()  ;
            end
            begin
              dma2mem[5][29].run()  ;
            end

            begin
              gen[5][30].run()  ;
            end
            begin
              drv[5][30].run()  ;
            end
            begin
              dma2mem[5][30].run()  ;
            end

            begin
              gen[5][31].run()  ;
            end
            begin
              drv[5][31].run()  ;
            end
            begin
              dma2mem[5][31].run()  ;
            end

            begin
              gen[6][0].run()  ;
            end
            begin
              drv[6][0].run()  ;
            end
            begin
              dma2mem[6][0].run()  ;
            end

            begin
              gen[6][1].run()  ;
            end
            begin
              drv[6][1].run()  ;
            end
            begin
              dma2mem[6][1].run()  ;
            end

            begin
              gen[6][2].run()  ;
            end
            begin
              drv[6][2].run()  ;
            end
            begin
              dma2mem[6][2].run()  ;
            end

            begin
              gen[6][3].run()  ;
            end
            begin
              drv[6][3].run()  ;
            end
            begin
              dma2mem[6][3].run()  ;
            end

            begin
              gen[6][4].run()  ;
            end
            begin
              drv[6][4].run()  ;
            end
            begin
              dma2mem[6][4].run()  ;
            end

            begin
              gen[6][5].run()  ;
            end
            begin
              drv[6][5].run()  ;
            end
            begin
              dma2mem[6][5].run()  ;
            end

            begin
              gen[6][6].run()  ;
            end
            begin
              drv[6][6].run()  ;
            end
            begin
              dma2mem[6][6].run()  ;
            end

            begin
              gen[6][7].run()  ;
            end
            begin
              drv[6][7].run()  ;
            end
            begin
              dma2mem[6][7].run()  ;
            end

            begin
              gen[6][8].run()  ;
            end
            begin
              drv[6][8].run()  ;
            end
            begin
              dma2mem[6][8].run()  ;
            end

            begin
              gen[6][9].run()  ;
            end
            begin
              drv[6][9].run()  ;
            end
            begin
              dma2mem[6][9].run()  ;
            end

            begin
              gen[6][10].run()  ;
            end
            begin
              drv[6][10].run()  ;
            end
            begin
              dma2mem[6][10].run()  ;
            end

            begin
              gen[6][11].run()  ;
            end
            begin
              drv[6][11].run()  ;
            end
            begin
              dma2mem[6][11].run()  ;
            end

            begin
              gen[6][12].run()  ;
            end
            begin
              drv[6][12].run()  ;
            end
            begin
              dma2mem[6][12].run()  ;
            end

            begin
              gen[6][13].run()  ;
            end
            begin
              drv[6][13].run()  ;
            end
            begin
              dma2mem[6][13].run()  ;
            end

            begin
              gen[6][14].run()  ;
            end
            begin
              drv[6][14].run()  ;
            end
            begin
              dma2mem[6][14].run()  ;
            end

            begin
              gen[6][15].run()  ;
            end
            begin
              drv[6][15].run()  ;
            end
            begin
              dma2mem[6][15].run()  ;
            end

            begin
              gen[6][16].run()  ;
            end
            begin
              drv[6][16].run()  ;
            end
            begin
              dma2mem[6][16].run()  ;
            end

            begin
              gen[6][17].run()  ;
            end
            begin
              drv[6][17].run()  ;
            end
            begin
              dma2mem[6][17].run()  ;
            end

            begin
              gen[6][18].run()  ;
            end
            begin
              drv[6][18].run()  ;
            end
            begin
              dma2mem[6][18].run()  ;
            end

            begin
              gen[6][19].run()  ;
            end
            begin
              drv[6][19].run()  ;
            end
            begin
              dma2mem[6][19].run()  ;
            end

            begin
              gen[6][20].run()  ;
            end
            begin
              drv[6][20].run()  ;
            end
            begin
              dma2mem[6][20].run()  ;
            end

            begin
              gen[6][21].run()  ;
            end
            begin
              drv[6][21].run()  ;
            end
            begin
              dma2mem[6][21].run()  ;
            end

            begin
              gen[6][22].run()  ;
            end
            begin
              drv[6][22].run()  ;
            end
            begin
              dma2mem[6][22].run()  ;
            end

            begin
              gen[6][23].run()  ;
            end
            begin
              drv[6][23].run()  ;
            end
            begin
              dma2mem[6][23].run()  ;
            end

            begin
              gen[6][24].run()  ;
            end
            begin
              drv[6][24].run()  ;
            end
            begin
              dma2mem[6][24].run()  ;
            end

            begin
              gen[6][25].run()  ;
            end
            begin
              drv[6][25].run()  ;
            end
            begin
              dma2mem[6][25].run()  ;
            end

            begin
              gen[6][26].run()  ;
            end
            begin
              drv[6][26].run()  ;
            end
            begin
              dma2mem[6][26].run()  ;
            end

            begin
              gen[6][27].run()  ;
            end
            begin
              drv[6][27].run()  ;
            end
            begin
              dma2mem[6][27].run()  ;
            end

            begin
              gen[6][28].run()  ;
            end
            begin
              drv[6][28].run()  ;
            end
            begin
              dma2mem[6][28].run()  ;
            end

            begin
              gen[6][29].run()  ;
            end
            begin
              drv[6][29].run()  ;
            end
            begin
              dma2mem[6][29].run()  ;
            end

            begin
              gen[6][30].run()  ;
            end
            begin
              drv[6][30].run()  ;
            end
            begin
              dma2mem[6][30].run()  ;
            end

            begin
              gen[6][31].run()  ;
            end
            begin
              drv[6][31].run()  ;
            end
            begin
              dma2mem[6][31].run()  ;
            end

            begin
              gen[7][0].run()  ;
            end
            begin
              drv[7][0].run()  ;
            end
            begin
              dma2mem[7][0].run()  ;
            end

            begin
              gen[7][1].run()  ;
            end
            begin
              drv[7][1].run()  ;
            end
            begin
              dma2mem[7][1].run()  ;
            end

            begin
              gen[7][2].run()  ;
            end
            begin
              drv[7][2].run()  ;
            end
            begin
              dma2mem[7][2].run()  ;
            end

            begin
              gen[7][3].run()  ;
            end
            begin
              drv[7][3].run()  ;
            end
            begin
              dma2mem[7][3].run()  ;
            end

            begin
              gen[7][4].run()  ;
            end
            begin
              drv[7][4].run()  ;
            end
            begin
              dma2mem[7][4].run()  ;
            end

            begin
              gen[7][5].run()  ;
            end
            begin
              drv[7][5].run()  ;
            end
            begin
              dma2mem[7][5].run()  ;
            end

            begin
              gen[7][6].run()  ;
            end
            begin
              drv[7][6].run()  ;
            end
            begin
              dma2mem[7][6].run()  ;
            end

            begin
              gen[7][7].run()  ;
            end
            begin
              drv[7][7].run()  ;
            end
            begin
              dma2mem[7][7].run()  ;
            end

            begin
              gen[7][8].run()  ;
            end
            begin
              drv[7][8].run()  ;
            end
            begin
              dma2mem[7][8].run()  ;
            end

            begin
              gen[7][9].run()  ;
            end
            begin
              drv[7][9].run()  ;
            end
            begin
              dma2mem[7][9].run()  ;
            end

            begin
              gen[7][10].run()  ;
            end
            begin
              drv[7][10].run()  ;
            end
            begin
              dma2mem[7][10].run()  ;
            end

            begin
              gen[7][11].run()  ;
            end
            begin
              drv[7][11].run()  ;
            end
            begin
              dma2mem[7][11].run()  ;
            end

            begin
              gen[7][12].run()  ;
            end
            begin
              drv[7][12].run()  ;
            end
            begin
              dma2mem[7][12].run()  ;
            end

            begin
              gen[7][13].run()  ;
            end
            begin
              drv[7][13].run()  ;
            end
            begin
              dma2mem[7][13].run()  ;
            end

            begin
              gen[7][14].run()  ;
            end
            begin
              drv[7][14].run()  ;
            end
            begin
              dma2mem[7][14].run()  ;
            end

            begin
              gen[7][15].run()  ;
            end
            begin
              drv[7][15].run()  ;
            end
            begin
              dma2mem[7][15].run()  ;
            end

            begin
              gen[7][16].run()  ;
            end
            begin
              drv[7][16].run()  ;
            end
            begin
              dma2mem[7][16].run()  ;
            end

            begin
              gen[7][17].run()  ;
            end
            begin
              drv[7][17].run()  ;
            end
            begin
              dma2mem[7][17].run()  ;
            end

            begin
              gen[7][18].run()  ;
            end
            begin
              drv[7][18].run()  ;
            end
            begin
              dma2mem[7][18].run()  ;
            end

            begin
              gen[7][19].run()  ;
            end
            begin
              drv[7][19].run()  ;
            end
            begin
              dma2mem[7][19].run()  ;
            end

            begin
              gen[7][20].run()  ;
            end
            begin
              drv[7][20].run()  ;
            end
            begin
              dma2mem[7][20].run()  ;
            end

            begin
              gen[7][21].run()  ;
            end
            begin
              drv[7][21].run()  ;
            end
            begin
              dma2mem[7][21].run()  ;
            end

            begin
              gen[7][22].run()  ;
            end
            begin
              drv[7][22].run()  ;
            end
            begin
              dma2mem[7][22].run()  ;
            end

            begin
              gen[7][23].run()  ;
            end
            begin
              drv[7][23].run()  ;
            end
            begin
              dma2mem[7][23].run()  ;
            end

            begin
              gen[7][24].run()  ;
            end
            begin
              drv[7][24].run()  ;
            end
            begin
              dma2mem[7][24].run()  ;
            end

            begin
              gen[7][25].run()  ;
            end
            begin
              drv[7][25].run()  ;
            end
            begin
              dma2mem[7][25].run()  ;
            end

            begin
              gen[7][26].run()  ;
            end
            begin
              drv[7][26].run()  ;
            end
            begin
              dma2mem[7][26].run()  ;
            end

            begin
              gen[7][27].run()  ;
            end
            begin
              drv[7][27].run()  ;
            end
            begin
              dma2mem[7][27].run()  ;
            end

            begin
              gen[7][28].run()  ;
            end
            begin
              drv[7][28].run()  ;
            end
            begin
              dma2mem[7][28].run()  ;
            end

            begin
              gen[7][29].run()  ;
            end
            begin
              drv[7][29].run()  ;
            end
            begin
              dma2mem[7][29].run()  ;
            end

            begin
              gen[7][30].run()  ;
            end
            begin
              drv[7][30].run()  ;
            end
            begin
              dma2mem[7][30].run()  ;
            end

            begin
              gen[7][31].run()  ;
            end
            begin
              drv[7][31].run()  ;
            end
            begin
              dma2mem[7][31].run()  ;
            end

            begin
              gen[8][0].run()  ;
            end
            begin
              drv[8][0].run()  ;
            end
            begin
              dma2mem[8][0].run()  ;
            end

            begin
              gen[8][1].run()  ;
            end
            begin
              drv[8][1].run()  ;
            end
            begin
              dma2mem[8][1].run()  ;
            end

            begin
              gen[8][2].run()  ;
            end
            begin
              drv[8][2].run()  ;
            end
            begin
              dma2mem[8][2].run()  ;
            end

            begin
              gen[8][3].run()  ;
            end
            begin
              drv[8][3].run()  ;
            end
            begin
              dma2mem[8][3].run()  ;
            end

            begin
              gen[8][4].run()  ;
            end
            begin
              drv[8][4].run()  ;
            end
            begin
              dma2mem[8][4].run()  ;
            end

            begin
              gen[8][5].run()  ;
            end
            begin
              drv[8][5].run()  ;
            end
            begin
              dma2mem[8][5].run()  ;
            end

            begin
              gen[8][6].run()  ;
            end
            begin
              drv[8][6].run()  ;
            end
            begin
              dma2mem[8][6].run()  ;
            end

            begin
              gen[8][7].run()  ;
            end
            begin
              drv[8][7].run()  ;
            end
            begin
              dma2mem[8][7].run()  ;
            end

            begin
              gen[8][8].run()  ;
            end
            begin
              drv[8][8].run()  ;
            end
            begin
              dma2mem[8][8].run()  ;
            end

            begin
              gen[8][9].run()  ;
            end
            begin
              drv[8][9].run()  ;
            end
            begin
              dma2mem[8][9].run()  ;
            end

            begin
              gen[8][10].run()  ;
            end
            begin
              drv[8][10].run()  ;
            end
            begin
              dma2mem[8][10].run()  ;
            end

            begin
              gen[8][11].run()  ;
            end
            begin
              drv[8][11].run()  ;
            end
            begin
              dma2mem[8][11].run()  ;
            end

            begin
              gen[8][12].run()  ;
            end
            begin
              drv[8][12].run()  ;
            end
            begin
              dma2mem[8][12].run()  ;
            end

            begin
              gen[8][13].run()  ;
            end
            begin
              drv[8][13].run()  ;
            end
            begin
              dma2mem[8][13].run()  ;
            end

            begin
              gen[8][14].run()  ;
            end
            begin
              drv[8][14].run()  ;
            end
            begin
              dma2mem[8][14].run()  ;
            end

            begin
              gen[8][15].run()  ;
            end
            begin
              drv[8][15].run()  ;
            end
            begin
              dma2mem[8][15].run()  ;
            end

            begin
              gen[8][16].run()  ;
            end
            begin
              drv[8][16].run()  ;
            end
            begin
              dma2mem[8][16].run()  ;
            end

            begin
              gen[8][17].run()  ;
            end
            begin
              drv[8][17].run()  ;
            end
            begin
              dma2mem[8][17].run()  ;
            end

            begin
              gen[8][18].run()  ;
            end
            begin
              drv[8][18].run()  ;
            end
            begin
              dma2mem[8][18].run()  ;
            end

            begin
              gen[8][19].run()  ;
            end
            begin
              drv[8][19].run()  ;
            end
            begin
              dma2mem[8][19].run()  ;
            end

            begin
              gen[8][20].run()  ;
            end
            begin
              drv[8][20].run()  ;
            end
            begin
              dma2mem[8][20].run()  ;
            end

            begin
              gen[8][21].run()  ;
            end
            begin
              drv[8][21].run()  ;
            end
            begin
              dma2mem[8][21].run()  ;
            end

            begin
              gen[8][22].run()  ;
            end
            begin
              drv[8][22].run()  ;
            end
            begin
              dma2mem[8][22].run()  ;
            end

            begin
              gen[8][23].run()  ;
            end
            begin
              drv[8][23].run()  ;
            end
            begin
              dma2mem[8][23].run()  ;
            end

            begin
              gen[8][24].run()  ;
            end
            begin
              drv[8][24].run()  ;
            end
            begin
              dma2mem[8][24].run()  ;
            end

            begin
              gen[8][25].run()  ;
            end
            begin
              drv[8][25].run()  ;
            end
            begin
              dma2mem[8][25].run()  ;
            end

            begin
              gen[8][26].run()  ;
            end
            begin
              drv[8][26].run()  ;
            end
            begin
              dma2mem[8][26].run()  ;
            end

            begin
              gen[8][27].run()  ;
            end
            begin
              drv[8][27].run()  ;
            end
            begin
              dma2mem[8][27].run()  ;
            end

            begin
              gen[8][28].run()  ;
            end
            begin
              drv[8][28].run()  ;
            end
            begin
              dma2mem[8][28].run()  ;
            end

            begin
              gen[8][29].run()  ;
            end
            begin
              drv[8][29].run()  ;
            end
            begin
              dma2mem[8][29].run()  ;
            end

            begin
              gen[8][30].run()  ;
            end
            begin
              drv[8][30].run()  ;
            end
            begin
              dma2mem[8][30].run()  ;
            end

            begin
              gen[8][31].run()  ;
            end
            begin
              drv[8][31].run()  ;
            end
            begin
              dma2mem[8][31].run()  ;
            end

            begin
              gen[9][0].run()  ;
            end
            begin
              drv[9][0].run()  ;
            end
            begin
              dma2mem[9][0].run()  ;
            end

            begin
              gen[9][1].run()  ;
            end
            begin
              drv[9][1].run()  ;
            end
            begin
              dma2mem[9][1].run()  ;
            end

            begin
              gen[9][2].run()  ;
            end
            begin
              drv[9][2].run()  ;
            end
            begin
              dma2mem[9][2].run()  ;
            end

            begin
              gen[9][3].run()  ;
            end
            begin
              drv[9][3].run()  ;
            end
            begin
              dma2mem[9][3].run()  ;
            end

            begin
              gen[9][4].run()  ;
            end
            begin
              drv[9][4].run()  ;
            end
            begin
              dma2mem[9][4].run()  ;
            end

            begin
              gen[9][5].run()  ;
            end
            begin
              drv[9][5].run()  ;
            end
            begin
              dma2mem[9][5].run()  ;
            end

            begin
              gen[9][6].run()  ;
            end
            begin
              drv[9][6].run()  ;
            end
            begin
              dma2mem[9][6].run()  ;
            end

            begin
              gen[9][7].run()  ;
            end
            begin
              drv[9][7].run()  ;
            end
            begin
              dma2mem[9][7].run()  ;
            end

            begin
              gen[9][8].run()  ;
            end
            begin
              drv[9][8].run()  ;
            end
            begin
              dma2mem[9][8].run()  ;
            end

            begin
              gen[9][9].run()  ;
            end
            begin
              drv[9][9].run()  ;
            end
            begin
              dma2mem[9][9].run()  ;
            end

            begin
              gen[9][10].run()  ;
            end
            begin
              drv[9][10].run()  ;
            end
            begin
              dma2mem[9][10].run()  ;
            end

            begin
              gen[9][11].run()  ;
            end
            begin
              drv[9][11].run()  ;
            end
            begin
              dma2mem[9][11].run()  ;
            end

            begin
              gen[9][12].run()  ;
            end
            begin
              drv[9][12].run()  ;
            end
            begin
              dma2mem[9][12].run()  ;
            end

            begin
              gen[9][13].run()  ;
            end
            begin
              drv[9][13].run()  ;
            end
            begin
              dma2mem[9][13].run()  ;
            end

            begin
              gen[9][14].run()  ;
            end
            begin
              drv[9][14].run()  ;
            end
            begin
              dma2mem[9][14].run()  ;
            end

            begin
              gen[9][15].run()  ;
            end
            begin
              drv[9][15].run()  ;
            end
            begin
              dma2mem[9][15].run()  ;
            end

            begin
              gen[9][16].run()  ;
            end
            begin
              drv[9][16].run()  ;
            end
            begin
              dma2mem[9][16].run()  ;
            end

            begin
              gen[9][17].run()  ;
            end
            begin
              drv[9][17].run()  ;
            end
            begin
              dma2mem[9][17].run()  ;
            end

            begin
              gen[9][18].run()  ;
            end
            begin
              drv[9][18].run()  ;
            end
            begin
              dma2mem[9][18].run()  ;
            end

            begin
              gen[9][19].run()  ;
            end
            begin
              drv[9][19].run()  ;
            end
            begin
              dma2mem[9][19].run()  ;
            end

            begin
              gen[9][20].run()  ;
            end
            begin
              drv[9][20].run()  ;
            end
            begin
              dma2mem[9][20].run()  ;
            end

            begin
              gen[9][21].run()  ;
            end
            begin
              drv[9][21].run()  ;
            end
            begin
              dma2mem[9][21].run()  ;
            end

            begin
              gen[9][22].run()  ;
            end
            begin
              drv[9][22].run()  ;
            end
            begin
              dma2mem[9][22].run()  ;
            end

            begin
              gen[9][23].run()  ;
            end
            begin
              drv[9][23].run()  ;
            end
            begin
              dma2mem[9][23].run()  ;
            end

            begin
              gen[9][24].run()  ;
            end
            begin
              drv[9][24].run()  ;
            end
            begin
              dma2mem[9][24].run()  ;
            end

            begin
              gen[9][25].run()  ;
            end
            begin
              drv[9][25].run()  ;
            end
            begin
              dma2mem[9][25].run()  ;
            end

            begin
              gen[9][26].run()  ;
            end
            begin
              drv[9][26].run()  ;
            end
            begin
              dma2mem[9][26].run()  ;
            end

            begin
              gen[9][27].run()  ;
            end
            begin
              drv[9][27].run()  ;
            end
            begin
              dma2mem[9][27].run()  ;
            end

            begin
              gen[9][28].run()  ;
            end
            begin
              drv[9][28].run()  ;
            end
            begin
              dma2mem[9][28].run()  ;
            end

            begin
              gen[9][29].run()  ;
            end
            begin
              drv[9][29].run()  ;
            end
            begin
              dma2mem[9][29].run()  ;
            end

            begin
              gen[9][30].run()  ;
            end
            begin
              drv[9][30].run()  ;
            end
            begin
              dma2mem[9][30].run()  ;
            end

            begin
              gen[9][31].run()  ;
            end
            begin
              drv[9][31].run()  ;
            end
            begin
              dma2mem[9][31].run()  ;
            end

            begin
              gen[10][0].run()  ;
            end
            begin
              drv[10][0].run()  ;
            end
            begin
              dma2mem[10][0].run()  ;
            end

            begin
              gen[10][1].run()  ;
            end
            begin
              drv[10][1].run()  ;
            end
            begin
              dma2mem[10][1].run()  ;
            end

            begin
              gen[10][2].run()  ;
            end
            begin
              drv[10][2].run()  ;
            end
            begin
              dma2mem[10][2].run()  ;
            end

            begin
              gen[10][3].run()  ;
            end
            begin
              drv[10][3].run()  ;
            end
            begin
              dma2mem[10][3].run()  ;
            end

            begin
              gen[10][4].run()  ;
            end
            begin
              drv[10][4].run()  ;
            end
            begin
              dma2mem[10][4].run()  ;
            end

            begin
              gen[10][5].run()  ;
            end
            begin
              drv[10][5].run()  ;
            end
            begin
              dma2mem[10][5].run()  ;
            end

            begin
              gen[10][6].run()  ;
            end
            begin
              drv[10][6].run()  ;
            end
            begin
              dma2mem[10][6].run()  ;
            end

            begin
              gen[10][7].run()  ;
            end
            begin
              drv[10][7].run()  ;
            end
            begin
              dma2mem[10][7].run()  ;
            end

            begin
              gen[10][8].run()  ;
            end
            begin
              drv[10][8].run()  ;
            end
            begin
              dma2mem[10][8].run()  ;
            end

            begin
              gen[10][9].run()  ;
            end
            begin
              drv[10][9].run()  ;
            end
            begin
              dma2mem[10][9].run()  ;
            end

            begin
              gen[10][10].run()  ;
            end
            begin
              drv[10][10].run()  ;
            end
            begin
              dma2mem[10][10].run()  ;
            end

            begin
              gen[10][11].run()  ;
            end
            begin
              drv[10][11].run()  ;
            end
            begin
              dma2mem[10][11].run()  ;
            end

            begin
              gen[10][12].run()  ;
            end
            begin
              drv[10][12].run()  ;
            end
            begin
              dma2mem[10][12].run()  ;
            end

            begin
              gen[10][13].run()  ;
            end
            begin
              drv[10][13].run()  ;
            end
            begin
              dma2mem[10][13].run()  ;
            end

            begin
              gen[10][14].run()  ;
            end
            begin
              drv[10][14].run()  ;
            end
            begin
              dma2mem[10][14].run()  ;
            end

            begin
              gen[10][15].run()  ;
            end
            begin
              drv[10][15].run()  ;
            end
            begin
              dma2mem[10][15].run()  ;
            end

            begin
              gen[10][16].run()  ;
            end
            begin
              drv[10][16].run()  ;
            end
            begin
              dma2mem[10][16].run()  ;
            end

            begin
              gen[10][17].run()  ;
            end
            begin
              drv[10][17].run()  ;
            end
            begin
              dma2mem[10][17].run()  ;
            end

            begin
              gen[10][18].run()  ;
            end
            begin
              drv[10][18].run()  ;
            end
            begin
              dma2mem[10][18].run()  ;
            end

            begin
              gen[10][19].run()  ;
            end
            begin
              drv[10][19].run()  ;
            end
            begin
              dma2mem[10][19].run()  ;
            end

            begin
              gen[10][20].run()  ;
            end
            begin
              drv[10][20].run()  ;
            end
            begin
              dma2mem[10][20].run()  ;
            end

            begin
              gen[10][21].run()  ;
            end
            begin
              drv[10][21].run()  ;
            end
            begin
              dma2mem[10][21].run()  ;
            end

            begin
              gen[10][22].run()  ;
            end
            begin
              drv[10][22].run()  ;
            end
            begin
              dma2mem[10][22].run()  ;
            end

            begin
              gen[10][23].run()  ;
            end
            begin
              drv[10][23].run()  ;
            end
            begin
              dma2mem[10][23].run()  ;
            end

            begin
              gen[10][24].run()  ;
            end
            begin
              drv[10][24].run()  ;
            end
            begin
              dma2mem[10][24].run()  ;
            end

            begin
              gen[10][25].run()  ;
            end
            begin
              drv[10][25].run()  ;
            end
            begin
              dma2mem[10][25].run()  ;
            end

            begin
              gen[10][26].run()  ;
            end
            begin
              drv[10][26].run()  ;
            end
            begin
              dma2mem[10][26].run()  ;
            end

            begin
              gen[10][27].run()  ;
            end
            begin
              drv[10][27].run()  ;
            end
            begin
              dma2mem[10][27].run()  ;
            end

            begin
              gen[10][28].run()  ;
            end
            begin
              drv[10][28].run()  ;
            end
            begin
              dma2mem[10][28].run()  ;
            end

            begin
              gen[10][29].run()  ;
            end
            begin
              drv[10][29].run()  ;
            end
            begin
              dma2mem[10][29].run()  ;
            end

            begin
              gen[10][30].run()  ;
            end
            begin
              drv[10][30].run()  ;
            end
            begin
              dma2mem[10][30].run()  ;
            end

            begin
              gen[10][31].run()  ;
            end
            begin
              drv[10][31].run()  ;
            end
            begin
              dma2mem[10][31].run()  ;
            end

            begin
              gen[11][0].run()  ;
            end
            begin
              drv[11][0].run()  ;
            end
            begin
              dma2mem[11][0].run()  ;
            end

            begin
              gen[11][1].run()  ;
            end
            begin
              drv[11][1].run()  ;
            end
            begin
              dma2mem[11][1].run()  ;
            end

            begin
              gen[11][2].run()  ;
            end
            begin
              drv[11][2].run()  ;
            end
            begin
              dma2mem[11][2].run()  ;
            end

            begin
              gen[11][3].run()  ;
            end
            begin
              drv[11][3].run()  ;
            end
            begin
              dma2mem[11][3].run()  ;
            end

            begin
              gen[11][4].run()  ;
            end
            begin
              drv[11][4].run()  ;
            end
            begin
              dma2mem[11][4].run()  ;
            end

            begin
              gen[11][5].run()  ;
            end
            begin
              drv[11][5].run()  ;
            end
            begin
              dma2mem[11][5].run()  ;
            end

            begin
              gen[11][6].run()  ;
            end
            begin
              drv[11][6].run()  ;
            end
            begin
              dma2mem[11][6].run()  ;
            end

            begin
              gen[11][7].run()  ;
            end
            begin
              drv[11][7].run()  ;
            end
            begin
              dma2mem[11][7].run()  ;
            end

            begin
              gen[11][8].run()  ;
            end
            begin
              drv[11][8].run()  ;
            end
            begin
              dma2mem[11][8].run()  ;
            end

            begin
              gen[11][9].run()  ;
            end
            begin
              drv[11][9].run()  ;
            end
            begin
              dma2mem[11][9].run()  ;
            end

            begin
              gen[11][10].run()  ;
            end
            begin
              drv[11][10].run()  ;
            end
            begin
              dma2mem[11][10].run()  ;
            end

            begin
              gen[11][11].run()  ;
            end
            begin
              drv[11][11].run()  ;
            end
            begin
              dma2mem[11][11].run()  ;
            end

            begin
              gen[11][12].run()  ;
            end
            begin
              drv[11][12].run()  ;
            end
            begin
              dma2mem[11][12].run()  ;
            end

            begin
              gen[11][13].run()  ;
            end
            begin
              drv[11][13].run()  ;
            end
            begin
              dma2mem[11][13].run()  ;
            end

            begin
              gen[11][14].run()  ;
            end
            begin
              drv[11][14].run()  ;
            end
            begin
              dma2mem[11][14].run()  ;
            end

            begin
              gen[11][15].run()  ;
            end
            begin
              drv[11][15].run()  ;
            end
            begin
              dma2mem[11][15].run()  ;
            end

            begin
              gen[11][16].run()  ;
            end
            begin
              drv[11][16].run()  ;
            end
            begin
              dma2mem[11][16].run()  ;
            end

            begin
              gen[11][17].run()  ;
            end
            begin
              drv[11][17].run()  ;
            end
            begin
              dma2mem[11][17].run()  ;
            end

            begin
              gen[11][18].run()  ;
            end
            begin
              drv[11][18].run()  ;
            end
            begin
              dma2mem[11][18].run()  ;
            end

            begin
              gen[11][19].run()  ;
            end
            begin
              drv[11][19].run()  ;
            end
            begin
              dma2mem[11][19].run()  ;
            end

            begin
              gen[11][20].run()  ;
            end
            begin
              drv[11][20].run()  ;
            end
            begin
              dma2mem[11][20].run()  ;
            end

            begin
              gen[11][21].run()  ;
            end
            begin
              drv[11][21].run()  ;
            end
            begin
              dma2mem[11][21].run()  ;
            end

            begin
              gen[11][22].run()  ;
            end
            begin
              drv[11][22].run()  ;
            end
            begin
              dma2mem[11][22].run()  ;
            end

            begin
              gen[11][23].run()  ;
            end
            begin
              drv[11][23].run()  ;
            end
            begin
              dma2mem[11][23].run()  ;
            end

            begin
              gen[11][24].run()  ;
            end
            begin
              drv[11][24].run()  ;
            end
            begin
              dma2mem[11][24].run()  ;
            end

            begin
              gen[11][25].run()  ;
            end
            begin
              drv[11][25].run()  ;
            end
            begin
              dma2mem[11][25].run()  ;
            end

            begin
              gen[11][26].run()  ;
            end
            begin
              drv[11][26].run()  ;
            end
            begin
              dma2mem[11][26].run()  ;
            end

            begin
              gen[11][27].run()  ;
            end
            begin
              drv[11][27].run()  ;
            end
            begin
              dma2mem[11][27].run()  ;
            end

            begin
              gen[11][28].run()  ;
            end
            begin
              drv[11][28].run()  ;
            end
            begin
              dma2mem[11][28].run()  ;
            end

            begin
              gen[11][29].run()  ;
            end
            begin
              drv[11][29].run()  ;
            end
            begin
              dma2mem[11][29].run()  ;
            end

            begin
              gen[11][30].run()  ;
            end
            begin
              drv[11][30].run()  ;
            end
            begin
              dma2mem[11][30].run()  ;
            end

            begin
              gen[11][31].run()  ;
            end
            begin
              drv[11][31].run()  ;
            end
            begin
              dma2mem[11][31].run()  ;
            end

            begin
              gen[12][0].run()  ;
            end
            begin
              drv[12][0].run()  ;
            end
            begin
              dma2mem[12][0].run()  ;
            end

            begin
              gen[12][1].run()  ;
            end
            begin
              drv[12][1].run()  ;
            end
            begin
              dma2mem[12][1].run()  ;
            end

            begin
              gen[12][2].run()  ;
            end
            begin
              drv[12][2].run()  ;
            end
            begin
              dma2mem[12][2].run()  ;
            end

            begin
              gen[12][3].run()  ;
            end
            begin
              drv[12][3].run()  ;
            end
            begin
              dma2mem[12][3].run()  ;
            end

            begin
              gen[12][4].run()  ;
            end
            begin
              drv[12][4].run()  ;
            end
            begin
              dma2mem[12][4].run()  ;
            end

            begin
              gen[12][5].run()  ;
            end
            begin
              drv[12][5].run()  ;
            end
            begin
              dma2mem[12][5].run()  ;
            end

            begin
              gen[12][6].run()  ;
            end
            begin
              drv[12][6].run()  ;
            end
            begin
              dma2mem[12][6].run()  ;
            end

            begin
              gen[12][7].run()  ;
            end
            begin
              drv[12][7].run()  ;
            end
            begin
              dma2mem[12][7].run()  ;
            end

            begin
              gen[12][8].run()  ;
            end
            begin
              drv[12][8].run()  ;
            end
            begin
              dma2mem[12][8].run()  ;
            end

            begin
              gen[12][9].run()  ;
            end
            begin
              drv[12][9].run()  ;
            end
            begin
              dma2mem[12][9].run()  ;
            end

            begin
              gen[12][10].run()  ;
            end
            begin
              drv[12][10].run()  ;
            end
            begin
              dma2mem[12][10].run()  ;
            end

            begin
              gen[12][11].run()  ;
            end
            begin
              drv[12][11].run()  ;
            end
            begin
              dma2mem[12][11].run()  ;
            end

            begin
              gen[12][12].run()  ;
            end
            begin
              drv[12][12].run()  ;
            end
            begin
              dma2mem[12][12].run()  ;
            end

            begin
              gen[12][13].run()  ;
            end
            begin
              drv[12][13].run()  ;
            end
            begin
              dma2mem[12][13].run()  ;
            end

            begin
              gen[12][14].run()  ;
            end
            begin
              drv[12][14].run()  ;
            end
            begin
              dma2mem[12][14].run()  ;
            end

            begin
              gen[12][15].run()  ;
            end
            begin
              drv[12][15].run()  ;
            end
            begin
              dma2mem[12][15].run()  ;
            end

            begin
              gen[12][16].run()  ;
            end
            begin
              drv[12][16].run()  ;
            end
            begin
              dma2mem[12][16].run()  ;
            end

            begin
              gen[12][17].run()  ;
            end
            begin
              drv[12][17].run()  ;
            end
            begin
              dma2mem[12][17].run()  ;
            end

            begin
              gen[12][18].run()  ;
            end
            begin
              drv[12][18].run()  ;
            end
            begin
              dma2mem[12][18].run()  ;
            end

            begin
              gen[12][19].run()  ;
            end
            begin
              drv[12][19].run()  ;
            end
            begin
              dma2mem[12][19].run()  ;
            end

            begin
              gen[12][20].run()  ;
            end
            begin
              drv[12][20].run()  ;
            end
            begin
              dma2mem[12][20].run()  ;
            end

            begin
              gen[12][21].run()  ;
            end
            begin
              drv[12][21].run()  ;
            end
            begin
              dma2mem[12][21].run()  ;
            end

            begin
              gen[12][22].run()  ;
            end
            begin
              drv[12][22].run()  ;
            end
            begin
              dma2mem[12][22].run()  ;
            end

            begin
              gen[12][23].run()  ;
            end
            begin
              drv[12][23].run()  ;
            end
            begin
              dma2mem[12][23].run()  ;
            end

            begin
              gen[12][24].run()  ;
            end
            begin
              drv[12][24].run()  ;
            end
            begin
              dma2mem[12][24].run()  ;
            end

            begin
              gen[12][25].run()  ;
            end
            begin
              drv[12][25].run()  ;
            end
            begin
              dma2mem[12][25].run()  ;
            end

            begin
              gen[12][26].run()  ;
            end
            begin
              drv[12][26].run()  ;
            end
            begin
              dma2mem[12][26].run()  ;
            end

            begin
              gen[12][27].run()  ;
            end
            begin
              drv[12][27].run()  ;
            end
            begin
              dma2mem[12][27].run()  ;
            end

            begin
              gen[12][28].run()  ;
            end
            begin
              drv[12][28].run()  ;
            end
            begin
              dma2mem[12][28].run()  ;
            end

            begin
              gen[12][29].run()  ;
            end
            begin
              drv[12][29].run()  ;
            end
            begin
              dma2mem[12][29].run()  ;
            end

            begin
              gen[12][30].run()  ;
            end
            begin
              drv[12][30].run()  ;
            end
            begin
              dma2mem[12][30].run()  ;
            end

            begin
              gen[12][31].run()  ;
            end
            begin
              drv[12][31].run()  ;
            end
            begin
              dma2mem[12][31].run()  ;
            end

            begin
              gen[13][0].run()  ;
            end
            begin
              drv[13][0].run()  ;
            end
            begin
              dma2mem[13][0].run()  ;
            end

            begin
              gen[13][1].run()  ;
            end
            begin
              drv[13][1].run()  ;
            end
            begin
              dma2mem[13][1].run()  ;
            end

            begin
              gen[13][2].run()  ;
            end
            begin
              drv[13][2].run()  ;
            end
            begin
              dma2mem[13][2].run()  ;
            end

            begin
              gen[13][3].run()  ;
            end
            begin
              drv[13][3].run()  ;
            end
            begin
              dma2mem[13][3].run()  ;
            end

            begin
              gen[13][4].run()  ;
            end
            begin
              drv[13][4].run()  ;
            end
            begin
              dma2mem[13][4].run()  ;
            end

            begin
              gen[13][5].run()  ;
            end
            begin
              drv[13][5].run()  ;
            end
            begin
              dma2mem[13][5].run()  ;
            end

            begin
              gen[13][6].run()  ;
            end
            begin
              drv[13][6].run()  ;
            end
            begin
              dma2mem[13][6].run()  ;
            end

            begin
              gen[13][7].run()  ;
            end
            begin
              drv[13][7].run()  ;
            end
            begin
              dma2mem[13][7].run()  ;
            end

            begin
              gen[13][8].run()  ;
            end
            begin
              drv[13][8].run()  ;
            end
            begin
              dma2mem[13][8].run()  ;
            end

            begin
              gen[13][9].run()  ;
            end
            begin
              drv[13][9].run()  ;
            end
            begin
              dma2mem[13][9].run()  ;
            end

            begin
              gen[13][10].run()  ;
            end
            begin
              drv[13][10].run()  ;
            end
            begin
              dma2mem[13][10].run()  ;
            end

            begin
              gen[13][11].run()  ;
            end
            begin
              drv[13][11].run()  ;
            end
            begin
              dma2mem[13][11].run()  ;
            end

            begin
              gen[13][12].run()  ;
            end
            begin
              drv[13][12].run()  ;
            end
            begin
              dma2mem[13][12].run()  ;
            end

            begin
              gen[13][13].run()  ;
            end
            begin
              drv[13][13].run()  ;
            end
            begin
              dma2mem[13][13].run()  ;
            end

            begin
              gen[13][14].run()  ;
            end
            begin
              drv[13][14].run()  ;
            end
            begin
              dma2mem[13][14].run()  ;
            end

            begin
              gen[13][15].run()  ;
            end
            begin
              drv[13][15].run()  ;
            end
            begin
              dma2mem[13][15].run()  ;
            end

            begin
              gen[13][16].run()  ;
            end
            begin
              drv[13][16].run()  ;
            end
            begin
              dma2mem[13][16].run()  ;
            end

            begin
              gen[13][17].run()  ;
            end
            begin
              drv[13][17].run()  ;
            end
            begin
              dma2mem[13][17].run()  ;
            end

            begin
              gen[13][18].run()  ;
            end
            begin
              drv[13][18].run()  ;
            end
            begin
              dma2mem[13][18].run()  ;
            end

            begin
              gen[13][19].run()  ;
            end
            begin
              drv[13][19].run()  ;
            end
            begin
              dma2mem[13][19].run()  ;
            end

            begin
              gen[13][20].run()  ;
            end
            begin
              drv[13][20].run()  ;
            end
            begin
              dma2mem[13][20].run()  ;
            end

            begin
              gen[13][21].run()  ;
            end
            begin
              drv[13][21].run()  ;
            end
            begin
              dma2mem[13][21].run()  ;
            end

            begin
              gen[13][22].run()  ;
            end
            begin
              drv[13][22].run()  ;
            end
            begin
              dma2mem[13][22].run()  ;
            end

            begin
              gen[13][23].run()  ;
            end
            begin
              drv[13][23].run()  ;
            end
            begin
              dma2mem[13][23].run()  ;
            end

            begin
              gen[13][24].run()  ;
            end
            begin
              drv[13][24].run()  ;
            end
            begin
              dma2mem[13][24].run()  ;
            end

            begin
              gen[13][25].run()  ;
            end
            begin
              drv[13][25].run()  ;
            end
            begin
              dma2mem[13][25].run()  ;
            end

            begin
              gen[13][26].run()  ;
            end
            begin
              drv[13][26].run()  ;
            end
            begin
              dma2mem[13][26].run()  ;
            end

            begin
              gen[13][27].run()  ;
            end
            begin
              drv[13][27].run()  ;
            end
            begin
              dma2mem[13][27].run()  ;
            end

            begin
              gen[13][28].run()  ;
            end
            begin
              drv[13][28].run()  ;
            end
            begin
              dma2mem[13][28].run()  ;
            end

            begin
              gen[13][29].run()  ;
            end
            begin
              drv[13][29].run()  ;
            end
            begin
              dma2mem[13][29].run()  ;
            end

            begin
              gen[13][30].run()  ;
            end
            begin
              drv[13][30].run()  ;
            end
            begin
              dma2mem[13][30].run()  ;
            end

            begin
              gen[13][31].run()  ;
            end
            begin
              drv[13][31].run()  ;
            end
            begin
              dma2mem[13][31].run()  ;
            end

            begin
              gen[14][0].run()  ;
            end
            begin
              drv[14][0].run()  ;
            end
            begin
              dma2mem[14][0].run()  ;
            end

            begin
              gen[14][1].run()  ;
            end
            begin
              drv[14][1].run()  ;
            end
            begin
              dma2mem[14][1].run()  ;
            end

            begin
              gen[14][2].run()  ;
            end
            begin
              drv[14][2].run()  ;
            end
            begin
              dma2mem[14][2].run()  ;
            end

            begin
              gen[14][3].run()  ;
            end
            begin
              drv[14][3].run()  ;
            end
            begin
              dma2mem[14][3].run()  ;
            end

            begin
              gen[14][4].run()  ;
            end
            begin
              drv[14][4].run()  ;
            end
            begin
              dma2mem[14][4].run()  ;
            end

            begin
              gen[14][5].run()  ;
            end
            begin
              drv[14][5].run()  ;
            end
            begin
              dma2mem[14][5].run()  ;
            end

            begin
              gen[14][6].run()  ;
            end
            begin
              drv[14][6].run()  ;
            end
            begin
              dma2mem[14][6].run()  ;
            end

            begin
              gen[14][7].run()  ;
            end
            begin
              drv[14][7].run()  ;
            end
            begin
              dma2mem[14][7].run()  ;
            end

            begin
              gen[14][8].run()  ;
            end
            begin
              drv[14][8].run()  ;
            end
            begin
              dma2mem[14][8].run()  ;
            end

            begin
              gen[14][9].run()  ;
            end
            begin
              drv[14][9].run()  ;
            end
            begin
              dma2mem[14][9].run()  ;
            end

            begin
              gen[14][10].run()  ;
            end
            begin
              drv[14][10].run()  ;
            end
            begin
              dma2mem[14][10].run()  ;
            end

            begin
              gen[14][11].run()  ;
            end
            begin
              drv[14][11].run()  ;
            end
            begin
              dma2mem[14][11].run()  ;
            end

            begin
              gen[14][12].run()  ;
            end
            begin
              drv[14][12].run()  ;
            end
            begin
              dma2mem[14][12].run()  ;
            end

            begin
              gen[14][13].run()  ;
            end
            begin
              drv[14][13].run()  ;
            end
            begin
              dma2mem[14][13].run()  ;
            end

            begin
              gen[14][14].run()  ;
            end
            begin
              drv[14][14].run()  ;
            end
            begin
              dma2mem[14][14].run()  ;
            end

            begin
              gen[14][15].run()  ;
            end
            begin
              drv[14][15].run()  ;
            end
            begin
              dma2mem[14][15].run()  ;
            end

            begin
              gen[14][16].run()  ;
            end
            begin
              drv[14][16].run()  ;
            end
            begin
              dma2mem[14][16].run()  ;
            end

            begin
              gen[14][17].run()  ;
            end
            begin
              drv[14][17].run()  ;
            end
            begin
              dma2mem[14][17].run()  ;
            end

            begin
              gen[14][18].run()  ;
            end
            begin
              drv[14][18].run()  ;
            end
            begin
              dma2mem[14][18].run()  ;
            end

            begin
              gen[14][19].run()  ;
            end
            begin
              drv[14][19].run()  ;
            end
            begin
              dma2mem[14][19].run()  ;
            end

            begin
              gen[14][20].run()  ;
            end
            begin
              drv[14][20].run()  ;
            end
            begin
              dma2mem[14][20].run()  ;
            end

            begin
              gen[14][21].run()  ;
            end
            begin
              drv[14][21].run()  ;
            end
            begin
              dma2mem[14][21].run()  ;
            end

            begin
              gen[14][22].run()  ;
            end
            begin
              drv[14][22].run()  ;
            end
            begin
              dma2mem[14][22].run()  ;
            end

            begin
              gen[14][23].run()  ;
            end
            begin
              drv[14][23].run()  ;
            end
            begin
              dma2mem[14][23].run()  ;
            end

            begin
              gen[14][24].run()  ;
            end
            begin
              drv[14][24].run()  ;
            end
            begin
              dma2mem[14][24].run()  ;
            end

            begin
              gen[14][25].run()  ;
            end
            begin
              drv[14][25].run()  ;
            end
            begin
              dma2mem[14][25].run()  ;
            end

            begin
              gen[14][26].run()  ;
            end
            begin
              drv[14][26].run()  ;
            end
            begin
              dma2mem[14][26].run()  ;
            end

            begin
              gen[14][27].run()  ;
            end
            begin
              drv[14][27].run()  ;
            end
            begin
              dma2mem[14][27].run()  ;
            end

            begin
              gen[14][28].run()  ;
            end
            begin
              drv[14][28].run()  ;
            end
            begin
              dma2mem[14][28].run()  ;
            end

            begin
              gen[14][29].run()  ;
            end
            begin
              drv[14][29].run()  ;
            end
            begin
              dma2mem[14][29].run()  ;
            end

            begin
              gen[14][30].run()  ;
            end
            begin
              drv[14][30].run()  ;
            end
            begin
              dma2mem[14][30].run()  ;
            end

            begin
              gen[14][31].run()  ;
            end
            begin
              drv[14][31].run()  ;
            end
            begin
              dma2mem[14][31].run()  ;
            end

            begin
              gen[15][0].run()  ;
            end
            begin
              drv[15][0].run()  ;
            end
            begin
              dma2mem[15][0].run()  ;
            end

            begin
              gen[15][1].run()  ;
            end
            begin
              drv[15][1].run()  ;
            end
            begin
              dma2mem[15][1].run()  ;
            end

            begin
              gen[15][2].run()  ;
            end
            begin
              drv[15][2].run()  ;
            end
            begin
              dma2mem[15][2].run()  ;
            end

            begin
              gen[15][3].run()  ;
            end
            begin
              drv[15][3].run()  ;
            end
            begin
              dma2mem[15][3].run()  ;
            end

            begin
              gen[15][4].run()  ;
            end
            begin
              drv[15][4].run()  ;
            end
            begin
              dma2mem[15][4].run()  ;
            end

            begin
              gen[15][5].run()  ;
            end
            begin
              drv[15][5].run()  ;
            end
            begin
              dma2mem[15][5].run()  ;
            end

            begin
              gen[15][6].run()  ;
            end
            begin
              drv[15][6].run()  ;
            end
            begin
              dma2mem[15][6].run()  ;
            end

            begin
              gen[15][7].run()  ;
            end
            begin
              drv[15][7].run()  ;
            end
            begin
              dma2mem[15][7].run()  ;
            end

            begin
              gen[15][8].run()  ;
            end
            begin
              drv[15][8].run()  ;
            end
            begin
              dma2mem[15][8].run()  ;
            end

            begin
              gen[15][9].run()  ;
            end
            begin
              drv[15][9].run()  ;
            end
            begin
              dma2mem[15][9].run()  ;
            end

            begin
              gen[15][10].run()  ;
            end
            begin
              drv[15][10].run()  ;
            end
            begin
              dma2mem[15][10].run()  ;
            end

            begin
              gen[15][11].run()  ;
            end
            begin
              drv[15][11].run()  ;
            end
            begin
              dma2mem[15][11].run()  ;
            end

            begin
              gen[15][12].run()  ;
            end
            begin
              drv[15][12].run()  ;
            end
            begin
              dma2mem[15][12].run()  ;
            end

            begin
              gen[15][13].run()  ;
            end
            begin
              drv[15][13].run()  ;
            end
            begin
              dma2mem[15][13].run()  ;
            end

            begin
              gen[15][14].run()  ;
            end
            begin
              drv[15][14].run()  ;
            end
            begin
              dma2mem[15][14].run()  ;
            end

            begin
              gen[15][15].run()  ;
            end
            begin
              drv[15][15].run()  ;
            end
            begin
              dma2mem[15][15].run()  ;
            end

            begin
              gen[15][16].run()  ;
            end
            begin
              drv[15][16].run()  ;
            end
            begin
              dma2mem[15][16].run()  ;
            end

            begin
              gen[15][17].run()  ;
            end
            begin
              drv[15][17].run()  ;
            end
            begin
              dma2mem[15][17].run()  ;
            end

            begin
              gen[15][18].run()  ;
            end
            begin
              drv[15][18].run()  ;
            end
            begin
              dma2mem[15][18].run()  ;
            end

            begin
              gen[15][19].run()  ;
            end
            begin
              drv[15][19].run()  ;
            end
            begin
              dma2mem[15][19].run()  ;
            end

            begin
              gen[15][20].run()  ;
            end
            begin
              drv[15][20].run()  ;
            end
            begin
              dma2mem[15][20].run()  ;
            end

            begin
              gen[15][21].run()  ;
            end
            begin
              drv[15][21].run()  ;
            end
            begin
              dma2mem[15][21].run()  ;
            end

            begin
              gen[15][22].run()  ;
            end
            begin
              drv[15][22].run()  ;
            end
            begin
              dma2mem[15][22].run()  ;
            end

            begin
              gen[15][23].run()  ;
            end
            begin
              drv[15][23].run()  ;
            end
            begin
              dma2mem[15][23].run()  ;
            end

            begin
              gen[15][24].run()  ;
            end
            begin
              drv[15][24].run()  ;
            end
            begin
              dma2mem[15][24].run()  ;
            end

            begin
              gen[15][25].run()  ;
            end
            begin
              drv[15][25].run()  ;
            end
            begin
              dma2mem[15][25].run()  ;
            end

            begin
              gen[15][26].run()  ;
            end
            begin
              drv[15][26].run()  ;
            end
            begin
              dma2mem[15][26].run()  ;
            end

            begin
              gen[15][27].run()  ;
            end
            begin
              drv[15][27].run()  ;
            end
            begin
              dma2mem[15][27].run()  ;
            end

            begin
              gen[15][28].run()  ;
            end
            begin
              drv[15][28].run()  ;
            end
            begin
              dma2mem[15][28].run()  ;
            end

            begin
              gen[15][29].run()  ;
            end
            begin
              drv[15][29].run()  ;
            end
            begin
              dma2mem[15][29].run()  ;
            end

            begin
              gen[15][30].run()  ;
            end
            begin
              drv[15][30].run()  ;
            end
            begin
              dma2mem[15][30].run()  ;
            end

            begin
              gen[15][31].run()  ;
            end
            begin
              drv[15][31].run()  ;
            end
            begin
              dma2mem[15][31].run()  ;
            end

            begin
              gen[16][0].run()  ;
            end
            begin
              drv[16][0].run()  ;
            end
            begin
              dma2mem[16][0].run()  ;
            end

            begin
              gen[16][1].run()  ;
            end
            begin
              drv[16][1].run()  ;
            end
            begin
              dma2mem[16][1].run()  ;
            end

            begin
              gen[16][2].run()  ;
            end
            begin
              drv[16][2].run()  ;
            end
            begin
              dma2mem[16][2].run()  ;
            end

            begin
              gen[16][3].run()  ;
            end
            begin
              drv[16][3].run()  ;
            end
            begin
              dma2mem[16][3].run()  ;
            end

            begin
              gen[16][4].run()  ;
            end
            begin
              drv[16][4].run()  ;
            end
            begin
              dma2mem[16][4].run()  ;
            end

            begin
              gen[16][5].run()  ;
            end
            begin
              drv[16][5].run()  ;
            end
            begin
              dma2mem[16][5].run()  ;
            end

            begin
              gen[16][6].run()  ;
            end
            begin
              drv[16][6].run()  ;
            end
            begin
              dma2mem[16][6].run()  ;
            end

            begin
              gen[16][7].run()  ;
            end
            begin
              drv[16][7].run()  ;
            end
            begin
              dma2mem[16][7].run()  ;
            end

            begin
              gen[16][8].run()  ;
            end
            begin
              drv[16][8].run()  ;
            end
            begin
              dma2mem[16][8].run()  ;
            end

            begin
              gen[16][9].run()  ;
            end
            begin
              drv[16][9].run()  ;
            end
            begin
              dma2mem[16][9].run()  ;
            end

            begin
              gen[16][10].run()  ;
            end
            begin
              drv[16][10].run()  ;
            end
            begin
              dma2mem[16][10].run()  ;
            end

            begin
              gen[16][11].run()  ;
            end
            begin
              drv[16][11].run()  ;
            end
            begin
              dma2mem[16][11].run()  ;
            end

            begin
              gen[16][12].run()  ;
            end
            begin
              drv[16][12].run()  ;
            end
            begin
              dma2mem[16][12].run()  ;
            end

            begin
              gen[16][13].run()  ;
            end
            begin
              drv[16][13].run()  ;
            end
            begin
              dma2mem[16][13].run()  ;
            end

            begin
              gen[16][14].run()  ;
            end
            begin
              drv[16][14].run()  ;
            end
            begin
              dma2mem[16][14].run()  ;
            end

            begin
              gen[16][15].run()  ;
            end
            begin
              drv[16][15].run()  ;
            end
            begin
              dma2mem[16][15].run()  ;
            end

            begin
              gen[16][16].run()  ;
            end
            begin
              drv[16][16].run()  ;
            end
            begin
              dma2mem[16][16].run()  ;
            end

            begin
              gen[16][17].run()  ;
            end
            begin
              drv[16][17].run()  ;
            end
            begin
              dma2mem[16][17].run()  ;
            end

            begin
              gen[16][18].run()  ;
            end
            begin
              drv[16][18].run()  ;
            end
            begin
              dma2mem[16][18].run()  ;
            end

            begin
              gen[16][19].run()  ;
            end
            begin
              drv[16][19].run()  ;
            end
            begin
              dma2mem[16][19].run()  ;
            end

            begin
              gen[16][20].run()  ;
            end
            begin
              drv[16][20].run()  ;
            end
            begin
              dma2mem[16][20].run()  ;
            end

            begin
              gen[16][21].run()  ;
            end
            begin
              drv[16][21].run()  ;
            end
            begin
              dma2mem[16][21].run()  ;
            end

            begin
              gen[16][22].run()  ;
            end
            begin
              drv[16][22].run()  ;
            end
            begin
              dma2mem[16][22].run()  ;
            end

            begin
              gen[16][23].run()  ;
            end
            begin
              drv[16][23].run()  ;
            end
            begin
              dma2mem[16][23].run()  ;
            end

            begin
              gen[16][24].run()  ;
            end
            begin
              drv[16][24].run()  ;
            end
            begin
              dma2mem[16][24].run()  ;
            end

            begin
              gen[16][25].run()  ;
            end
            begin
              drv[16][25].run()  ;
            end
            begin
              dma2mem[16][25].run()  ;
            end

            begin
              gen[16][26].run()  ;
            end
            begin
              drv[16][26].run()  ;
            end
            begin
              dma2mem[16][26].run()  ;
            end

            begin
              gen[16][27].run()  ;
            end
            begin
              drv[16][27].run()  ;
            end
            begin
              dma2mem[16][27].run()  ;
            end

            begin
              gen[16][28].run()  ;
            end
            begin
              drv[16][28].run()  ;
            end
            begin
              dma2mem[16][28].run()  ;
            end

            begin
              gen[16][29].run()  ;
            end
            begin
              drv[16][29].run()  ;
            end
            begin
              dma2mem[16][29].run()  ;
            end

            begin
              gen[16][30].run()  ;
            end
            begin
              drv[16][30].run()  ;
            end
            begin
              dma2mem[16][30].run()  ;
            end

            begin
              gen[16][31].run()  ;
            end
            begin
              drv[16][31].run()  ;
            end
            begin
              dma2mem[16][31].run()  ;
            end

            begin
              gen[17][0].run()  ;
            end
            begin
              drv[17][0].run()  ;
            end
            begin
              dma2mem[17][0].run()  ;
            end

            begin
              gen[17][1].run()  ;
            end
            begin
              drv[17][1].run()  ;
            end
            begin
              dma2mem[17][1].run()  ;
            end

            begin
              gen[17][2].run()  ;
            end
            begin
              drv[17][2].run()  ;
            end
            begin
              dma2mem[17][2].run()  ;
            end

            begin
              gen[17][3].run()  ;
            end
            begin
              drv[17][3].run()  ;
            end
            begin
              dma2mem[17][3].run()  ;
            end

            begin
              gen[17][4].run()  ;
            end
            begin
              drv[17][4].run()  ;
            end
            begin
              dma2mem[17][4].run()  ;
            end

            begin
              gen[17][5].run()  ;
            end
            begin
              drv[17][5].run()  ;
            end
            begin
              dma2mem[17][5].run()  ;
            end

            begin
              gen[17][6].run()  ;
            end
            begin
              drv[17][6].run()  ;
            end
            begin
              dma2mem[17][6].run()  ;
            end

            begin
              gen[17][7].run()  ;
            end
            begin
              drv[17][7].run()  ;
            end
            begin
              dma2mem[17][7].run()  ;
            end

            begin
              gen[17][8].run()  ;
            end
            begin
              drv[17][8].run()  ;
            end
            begin
              dma2mem[17][8].run()  ;
            end

            begin
              gen[17][9].run()  ;
            end
            begin
              drv[17][9].run()  ;
            end
            begin
              dma2mem[17][9].run()  ;
            end

            begin
              gen[17][10].run()  ;
            end
            begin
              drv[17][10].run()  ;
            end
            begin
              dma2mem[17][10].run()  ;
            end

            begin
              gen[17][11].run()  ;
            end
            begin
              drv[17][11].run()  ;
            end
            begin
              dma2mem[17][11].run()  ;
            end

            begin
              gen[17][12].run()  ;
            end
            begin
              drv[17][12].run()  ;
            end
            begin
              dma2mem[17][12].run()  ;
            end

            begin
              gen[17][13].run()  ;
            end
            begin
              drv[17][13].run()  ;
            end
            begin
              dma2mem[17][13].run()  ;
            end

            begin
              gen[17][14].run()  ;
            end
            begin
              drv[17][14].run()  ;
            end
            begin
              dma2mem[17][14].run()  ;
            end

            begin
              gen[17][15].run()  ;
            end
            begin
              drv[17][15].run()  ;
            end
            begin
              dma2mem[17][15].run()  ;
            end

            begin
              gen[17][16].run()  ;
            end
            begin
              drv[17][16].run()  ;
            end
            begin
              dma2mem[17][16].run()  ;
            end

            begin
              gen[17][17].run()  ;
            end
            begin
              drv[17][17].run()  ;
            end
            begin
              dma2mem[17][17].run()  ;
            end

            begin
              gen[17][18].run()  ;
            end
            begin
              drv[17][18].run()  ;
            end
            begin
              dma2mem[17][18].run()  ;
            end

            begin
              gen[17][19].run()  ;
            end
            begin
              drv[17][19].run()  ;
            end
            begin
              dma2mem[17][19].run()  ;
            end

            begin
              gen[17][20].run()  ;
            end
            begin
              drv[17][20].run()  ;
            end
            begin
              dma2mem[17][20].run()  ;
            end

            begin
              gen[17][21].run()  ;
            end
            begin
              drv[17][21].run()  ;
            end
            begin
              dma2mem[17][21].run()  ;
            end

            begin
              gen[17][22].run()  ;
            end
            begin
              drv[17][22].run()  ;
            end
            begin
              dma2mem[17][22].run()  ;
            end

            begin
              gen[17][23].run()  ;
            end
            begin
              drv[17][23].run()  ;
            end
            begin
              dma2mem[17][23].run()  ;
            end

            begin
              gen[17][24].run()  ;
            end
            begin
              drv[17][24].run()  ;
            end
            begin
              dma2mem[17][24].run()  ;
            end

            begin
              gen[17][25].run()  ;
            end
            begin
              drv[17][25].run()  ;
            end
            begin
              dma2mem[17][25].run()  ;
            end

            begin
              gen[17][26].run()  ;
            end
            begin
              drv[17][26].run()  ;
            end
            begin
              dma2mem[17][26].run()  ;
            end

            begin
              gen[17][27].run()  ;
            end
            begin
              drv[17][27].run()  ;
            end
            begin
              dma2mem[17][27].run()  ;
            end

            begin
              gen[17][28].run()  ;
            end
            begin
              drv[17][28].run()  ;
            end
            begin
              dma2mem[17][28].run()  ;
            end

            begin
              gen[17][29].run()  ;
            end
            begin
              drv[17][29].run()  ;
            end
            begin
              dma2mem[17][29].run()  ;
            end

            begin
              gen[17][30].run()  ;
            end
            begin
              drv[17][30].run()  ;
            end
            begin
              dma2mem[17][30].run()  ;
            end

            begin
              gen[17][31].run()  ;
            end
            begin
              drv[17][31].run()  ;
            end
            begin
              dma2mem[17][31].run()  ;
            end

            begin
              gen[18][0].run()  ;
            end
            begin
              drv[18][0].run()  ;
            end
            begin
              dma2mem[18][0].run()  ;
            end

            begin
              gen[18][1].run()  ;
            end
            begin
              drv[18][1].run()  ;
            end
            begin
              dma2mem[18][1].run()  ;
            end

            begin
              gen[18][2].run()  ;
            end
            begin
              drv[18][2].run()  ;
            end
            begin
              dma2mem[18][2].run()  ;
            end

            begin
              gen[18][3].run()  ;
            end
            begin
              drv[18][3].run()  ;
            end
            begin
              dma2mem[18][3].run()  ;
            end

            begin
              gen[18][4].run()  ;
            end
            begin
              drv[18][4].run()  ;
            end
            begin
              dma2mem[18][4].run()  ;
            end

            begin
              gen[18][5].run()  ;
            end
            begin
              drv[18][5].run()  ;
            end
            begin
              dma2mem[18][5].run()  ;
            end

            begin
              gen[18][6].run()  ;
            end
            begin
              drv[18][6].run()  ;
            end
            begin
              dma2mem[18][6].run()  ;
            end

            begin
              gen[18][7].run()  ;
            end
            begin
              drv[18][7].run()  ;
            end
            begin
              dma2mem[18][7].run()  ;
            end

            begin
              gen[18][8].run()  ;
            end
            begin
              drv[18][8].run()  ;
            end
            begin
              dma2mem[18][8].run()  ;
            end

            begin
              gen[18][9].run()  ;
            end
            begin
              drv[18][9].run()  ;
            end
            begin
              dma2mem[18][9].run()  ;
            end

            begin
              gen[18][10].run()  ;
            end
            begin
              drv[18][10].run()  ;
            end
            begin
              dma2mem[18][10].run()  ;
            end

            begin
              gen[18][11].run()  ;
            end
            begin
              drv[18][11].run()  ;
            end
            begin
              dma2mem[18][11].run()  ;
            end

            begin
              gen[18][12].run()  ;
            end
            begin
              drv[18][12].run()  ;
            end
            begin
              dma2mem[18][12].run()  ;
            end

            begin
              gen[18][13].run()  ;
            end
            begin
              drv[18][13].run()  ;
            end
            begin
              dma2mem[18][13].run()  ;
            end

            begin
              gen[18][14].run()  ;
            end
            begin
              drv[18][14].run()  ;
            end
            begin
              dma2mem[18][14].run()  ;
            end

            begin
              gen[18][15].run()  ;
            end
            begin
              drv[18][15].run()  ;
            end
            begin
              dma2mem[18][15].run()  ;
            end

            begin
              gen[18][16].run()  ;
            end
            begin
              drv[18][16].run()  ;
            end
            begin
              dma2mem[18][16].run()  ;
            end

            begin
              gen[18][17].run()  ;
            end
            begin
              drv[18][17].run()  ;
            end
            begin
              dma2mem[18][17].run()  ;
            end

            begin
              gen[18][18].run()  ;
            end
            begin
              drv[18][18].run()  ;
            end
            begin
              dma2mem[18][18].run()  ;
            end

            begin
              gen[18][19].run()  ;
            end
            begin
              drv[18][19].run()  ;
            end
            begin
              dma2mem[18][19].run()  ;
            end

            begin
              gen[18][20].run()  ;
            end
            begin
              drv[18][20].run()  ;
            end
            begin
              dma2mem[18][20].run()  ;
            end

            begin
              gen[18][21].run()  ;
            end
            begin
              drv[18][21].run()  ;
            end
            begin
              dma2mem[18][21].run()  ;
            end

            begin
              gen[18][22].run()  ;
            end
            begin
              drv[18][22].run()  ;
            end
            begin
              dma2mem[18][22].run()  ;
            end

            begin
              gen[18][23].run()  ;
            end
            begin
              drv[18][23].run()  ;
            end
            begin
              dma2mem[18][23].run()  ;
            end

            begin
              gen[18][24].run()  ;
            end
            begin
              drv[18][24].run()  ;
            end
            begin
              dma2mem[18][24].run()  ;
            end

            begin
              gen[18][25].run()  ;
            end
            begin
              drv[18][25].run()  ;
            end
            begin
              dma2mem[18][25].run()  ;
            end

            begin
              gen[18][26].run()  ;
            end
            begin
              drv[18][26].run()  ;
            end
            begin
              dma2mem[18][26].run()  ;
            end

            begin
              gen[18][27].run()  ;
            end
            begin
              drv[18][27].run()  ;
            end
            begin
              dma2mem[18][27].run()  ;
            end

            begin
              gen[18][28].run()  ;
            end
            begin
              drv[18][28].run()  ;
            end
            begin
              dma2mem[18][28].run()  ;
            end

            begin
              gen[18][29].run()  ;
            end
            begin
              drv[18][29].run()  ;
            end
            begin
              dma2mem[18][29].run()  ;
            end

            begin
              gen[18][30].run()  ;
            end
            begin
              drv[18][30].run()  ;
            end
            begin
              dma2mem[18][30].run()  ;
            end

            begin
              gen[18][31].run()  ;
            end
            begin
              drv[18][31].run()  ;
            end
            begin
              dma2mem[18][31].run()  ;
            end

            begin
              gen[19][0].run()  ;
            end
            begin
              drv[19][0].run()  ;
            end
            begin
              dma2mem[19][0].run()  ;
            end

            begin
              gen[19][1].run()  ;
            end
            begin
              drv[19][1].run()  ;
            end
            begin
              dma2mem[19][1].run()  ;
            end

            begin
              gen[19][2].run()  ;
            end
            begin
              drv[19][2].run()  ;
            end
            begin
              dma2mem[19][2].run()  ;
            end

            begin
              gen[19][3].run()  ;
            end
            begin
              drv[19][3].run()  ;
            end
            begin
              dma2mem[19][3].run()  ;
            end

            begin
              gen[19][4].run()  ;
            end
            begin
              drv[19][4].run()  ;
            end
            begin
              dma2mem[19][4].run()  ;
            end

            begin
              gen[19][5].run()  ;
            end
            begin
              drv[19][5].run()  ;
            end
            begin
              dma2mem[19][5].run()  ;
            end

            begin
              gen[19][6].run()  ;
            end
            begin
              drv[19][6].run()  ;
            end
            begin
              dma2mem[19][6].run()  ;
            end

            begin
              gen[19][7].run()  ;
            end
            begin
              drv[19][7].run()  ;
            end
            begin
              dma2mem[19][7].run()  ;
            end

            begin
              gen[19][8].run()  ;
            end
            begin
              drv[19][8].run()  ;
            end
            begin
              dma2mem[19][8].run()  ;
            end

            begin
              gen[19][9].run()  ;
            end
            begin
              drv[19][9].run()  ;
            end
            begin
              dma2mem[19][9].run()  ;
            end

            begin
              gen[19][10].run()  ;
            end
            begin
              drv[19][10].run()  ;
            end
            begin
              dma2mem[19][10].run()  ;
            end

            begin
              gen[19][11].run()  ;
            end
            begin
              drv[19][11].run()  ;
            end
            begin
              dma2mem[19][11].run()  ;
            end

            begin
              gen[19][12].run()  ;
            end
            begin
              drv[19][12].run()  ;
            end
            begin
              dma2mem[19][12].run()  ;
            end

            begin
              gen[19][13].run()  ;
            end
            begin
              drv[19][13].run()  ;
            end
            begin
              dma2mem[19][13].run()  ;
            end

            begin
              gen[19][14].run()  ;
            end
            begin
              drv[19][14].run()  ;
            end
            begin
              dma2mem[19][14].run()  ;
            end

            begin
              gen[19][15].run()  ;
            end
            begin
              drv[19][15].run()  ;
            end
            begin
              dma2mem[19][15].run()  ;
            end

            begin
              gen[19][16].run()  ;
            end
            begin
              drv[19][16].run()  ;
            end
            begin
              dma2mem[19][16].run()  ;
            end

            begin
              gen[19][17].run()  ;
            end
            begin
              drv[19][17].run()  ;
            end
            begin
              dma2mem[19][17].run()  ;
            end

            begin
              gen[19][18].run()  ;
            end
            begin
              drv[19][18].run()  ;
            end
            begin
              dma2mem[19][18].run()  ;
            end

            begin
              gen[19][19].run()  ;
            end
            begin
              drv[19][19].run()  ;
            end
            begin
              dma2mem[19][19].run()  ;
            end

            begin
              gen[19][20].run()  ;
            end
            begin
              drv[19][20].run()  ;
            end
            begin
              dma2mem[19][20].run()  ;
            end

            begin
              gen[19][21].run()  ;
            end
            begin
              drv[19][21].run()  ;
            end
            begin
              dma2mem[19][21].run()  ;
            end

            begin
              gen[19][22].run()  ;
            end
            begin
              drv[19][22].run()  ;
            end
            begin
              dma2mem[19][22].run()  ;
            end

            begin
              gen[19][23].run()  ;
            end
            begin
              drv[19][23].run()  ;
            end
            begin
              dma2mem[19][23].run()  ;
            end

            begin
              gen[19][24].run()  ;
            end
            begin
              drv[19][24].run()  ;
            end
            begin
              dma2mem[19][24].run()  ;
            end

            begin
              gen[19][25].run()  ;
            end
            begin
              drv[19][25].run()  ;
            end
            begin
              dma2mem[19][25].run()  ;
            end

            begin
              gen[19][26].run()  ;
            end
            begin
              drv[19][26].run()  ;
            end
            begin
              dma2mem[19][26].run()  ;
            end

            begin
              gen[19][27].run()  ;
            end
            begin
              drv[19][27].run()  ;
            end
            begin
              dma2mem[19][27].run()  ;
            end

            begin
              gen[19][28].run()  ;
            end
            begin
              drv[19][28].run()  ;
            end
            begin
              dma2mem[19][28].run()  ;
            end

            begin
              gen[19][29].run()  ;
            end
            begin
              drv[19][29].run()  ;
            end
            begin
              dma2mem[19][29].run()  ;
            end

            begin
              gen[19][30].run()  ;
            end
            begin
              drv[19][30].run()  ;
            end
            begin
              dma2mem[19][30].run()  ;
            end

            begin
              gen[19][31].run()  ;
            end
            begin
              drv[19][31].run()  ;
            end
            begin
              dma2mem[19][31].run()  ;
            end

            begin
              gen[20][0].run()  ;
            end
            begin
              drv[20][0].run()  ;
            end
            begin
              dma2mem[20][0].run()  ;
            end

            begin
              gen[20][1].run()  ;
            end
            begin
              drv[20][1].run()  ;
            end
            begin
              dma2mem[20][1].run()  ;
            end

            begin
              gen[20][2].run()  ;
            end
            begin
              drv[20][2].run()  ;
            end
            begin
              dma2mem[20][2].run()  ;
            end

            begin
              gen[20][3].run()  ;
            end
            begin
              drv[20][3].run()  ;
            end
            begin
              dma2mem[20][3].run()  ;
            end

            begin
              gen[20][4].run()  ;
            end
            begin
              drv[20][4].run()  ;
            end
            begin
              dma2mem[20][4].run()  ;
            end

            begin
              gen[20][5].run()  ;
            end
            begin
              drv[20][5].run()  ;
            end
            begin
              dma2mem[20][5].run()  ;
            end

            begin
              gen[20][6].run()  ;
            end
            begin
              drv[20][6].run()  ;
            end
            begin
              dma2mem[20][6].run()  ;
            end

            begin
              gen[20][7].run()  ;
            end
            begin
              drv[20][7].run()  ;
            end
            begin
              dma2mem[20][7].run()  ;
            end

            begin
              gen[20][8].run()  ;
            end
            begin
              drv[20][8].run()  ;
            end
            begin
              dma2mem[20][8].run()  ;
            end

            begin
              gen[20][9].run()  ;
            end
            begin
              drv[20][9].run()  ;
            end
            begin
              dma2mem[20][9].run()  ;
            end

            begin
              gen[20][10].run()  ;
            end
            begin
              drv[20][10].run()  ;
            end
            begin
              dma2mem[20][10].run()  ;
            end

            begin
              gen[20][11].run()  ;
            end
            begin
              drv[20][11].run()  ;
            end
            begin
              dma2mem[20][11].run()  ;
            end

            begin
              gen[20][12].run()  ;
            end
            begin
              drv[20][12].run()  ;
            end
            begin
              dma2mem[20][12].run()  ;
            end

            begin
              gen[20][13].run()  ;
            end
            begin
              drv[20][13].run()  ;
            end
            begin
              dma2mem[20][13].run()  ;
            end

            begin
              gen[20][14].run()  ;
            end
            begin
              drv[20][14].run()  ;
            end
            begin
              dma2mem[20][14].run()  ;
            end

            begin
              gen[20][15].run()  ;
            end
            begin
              drv[20][15].run()  ;
            end
            begin
              dma2mem[20][15].run()  ;
            end

            begin
              gen[20][16].run()  ;
            end
            begin
              drv[20][16].run()  ;
            end
            begin
              dma2mem[20][16].run()  ;
            end

            begin
              gen[20][17].run()  ;
            end
            begin
              drv[20][17].run()  ;
            end
            begin
              dma2mem[20][17].run()  ;
            end

            begin
              gen[20][18].run()  ;
            end
            begin
              drv[20][18].run()  ;
            end
            begin
              dma2mem[20][18].run()  ;
            end

            begin
              gen[20][19].run()  ;
            end
            begin
              drv[20][19].run()  ;
            end
            begin
              dma2mem[20][19].run()  ;
            end

            begin
              gen[20][20].run()  ;
            end
            begin
              drv[20][20].run()  ;
            end
            begin
              dma2mem[20][20].run()  ;
            end

            begin
              gen[20][21].run()  ;
            end
            begin
              drv[20][21].run()  ;
            end
            begin
              dma2mem[20][21].run()  ;
            end

            begin
              gen[20][22].run()  ;
            end
            begin
              drv[20][22].run()  ;
            end
            begin
              dma2mem[20][22].run()  ;
            end

            begin
              gen[20][23].run()  ;
            end
            begin
              drv[20][23].run()  ;
            end
            begin
              dma2mem[20][23].run()  ;
            end

            begin
              gen[20][24].run()  ;
            end
            begin
              drv[20][24].run()  ;
            end
            begin
              dma2mem[20][24].run()  ;
            end

            begin
              gen[20][25].run()  ;
            end
            begin
              drv[20][25].run()  ;
            end
            begin
              dma2mem[20][25].run()  ;
            end

            begin
              gen[20][26].run()  ;
            end
            begin
              drv[20][26].run()  ;
            end
            begin
              dma2mem[20][26].run()  ;
            end

            begin
              gen[20][27].run()  ;
            end
            begin
              drv[20][27].run()  ;
            end
            begin
              dma2mem[20][27].run()  ;
            end

            begin
              gen[20][28].run()  ;
            end
            begin
              drv[20][28].run()  ;
            end
            begin
              dma2mem[20][28].run()  ;
            end

            begin
              gen[20][29].run()  ;
            end
            begin
              drv[20][29].run()  ;
            end
            begin
              dma2mem[20][29].run()  ;
            end

            begin
              gen[20][30].run()  ;
            end
            begin
              drv[20][30].run()  ;
            end
            begin
              dma2mem[20][30].run()  ;
            end

            begin
              gen[20][31].run()  ;
            end
            begin
              drv[20][31].run()  ;
            end
            begin
              dma2mem[20][31].run()  ;
            end

            begin
              gen[21][0].run()  ;
            end
            begin
              drv[21][0].run()  ;
            end
            begin
              dma2mem[21][0].run()  ;
            end

            begin
              gen[21][1].run()  ;
            end
            begin
              drv[21][1].run()  ;
            end
            begin
              dma2mem[21][1].run()  ;
            end

            begin
              gen[21][2].run()  ;
            end
            begin
              drv[21][2].run()  ;
            end
            begin
              dma2mem[21][2].run()  ;
            end

            begin
              gen[21][3].run()  ;
            end
            begin
              drv[21][3].run()  ;
            end
            begin
              dma2mem[21][3].run()  ;
            end

            begin
              gen[21][4].run()  ;
            end
            begin
              drv[21][4].run()  ;
            end
            begin
              dma2mem[21][4].run()  ;
            end

            begin
              gen[21][5].run()  ;
            end
            begin
              drv[21][5].run()  ;
            end
            begin
              dma2mem[21][5].run()  ;
            end

            begin
              gen[21][6].run()  ;
            end
            begin
              drv[21][6].run()  ;
            end
            begin
              dma2mem[21][6].run()  ;
            end

            begin
              gen[21][7].run()  ;
            end
            begin
              drv[21][7].run()  ;
            end
            begin
              dma2mem[21][7].run()  ;
            end

            begin
              gen[21][8].run()  ;
            end
            begin
              drv[21][8].run()  ;
            end
            begin
              dma2mem[21][8].run()  ;
            end

            begin
              gen[21][9].run()  ;
            end
            begin
              drv[21][9].run()  ;
            end
            begin
              dma2mem[21][9].run()  ;
            end

            begin
              gen[21][10].run()  ;
            end
            begin
              drv[21][10].run()  ;
            end
            begin
              dma2mem[21][10].run()  ;
            end

            begin
              gen[21][11].run()  ;
            end
            begin
              drv[21][11].run()  ;
            end
            begin
              dma2mem[21][11].run()  ;
            end

            begin
              gen[21][12].run()  ;
            end
            begin
              drv[21][12].run()  ;
            end
            begin
              dma2mem[21][12].run()  ;
            end

            begin
              gen[21][13].run()  ;
            end
            begin
              drv[21][13].run()  ;
            end
            begin
              dma2mem[21][13].run()  ;
            end

            begin
              gen[21][14].run()  ;
            end
            begin
              drv[21][14].run()  ;
            end
            begin
              dma2mem[21][14].run()  ;
            end

            begin
              gen[21][15].run()  ;
            end
            begin
              drv[21][15].run()  ;
            end
            begin
              dma2mem[21][15].run()  ;
            end

            begin
              gen[21][16].run()  ;
            end
            begin
              drv[21][16].run()  ;
            end
            begin
              dma2mem[21][16].run()  ;
            end

            begin
              gen[21][17].run()  ;
            end
            begin
              drv[21][17].run()  ;
            end
            begin
              dma2mem[21][17].run()  ;
            end

            begin
              gen[21][18].run()  ;
            end
            begin
              drv[21][18].run()  ;
            end
            begin
              dma2mem[21][18].run()  ;
            end

            begin
              gen[21][19].run()  ;
            end
            begin
              drv[21][19].run()  ;
            end
            begin
              dma2mem[21][19].run()  ;
            end

            begin
              gen[21][20].run()  ;
            end
            begin
              drv[21][20].run()  ;
            end
            begin
              dma2mem[21][20].run()  ;
            end

            begin
              gen[21][21].run()  ;
            end
            begin
              drv[21][21].run()  ;
            end
            begin
              dma2mem[21][21].run()  ;
            end

            begin
              gen[21][22].run()  ;
            end
            begin
              drv[21][22].run()  ;
            end
            begin
              dma2mem[21][22].run()  ;
            end

            begin
              gen[21][23].run()  ;
            end
            begin
              drv[21][23].run()  ;
            end
            begin
              dma2mem[21][23].run()  ;
            end

            begin
              gen[21][24].run()  ;
            end
            begin
              drv[21][24].run()  ;
            end
            begin
              dma2mem[21][24].run()  ;
            end

            begin
              gen[21][25].run()  ;
            end
            begin
              drv[21][25].run()  ;
            end
            begin
              dma2mem[21][25].run()  ;
            end

            begin
              gen[21][26].run()  ;
            end
            begin
              drv[21][26].run()  ;
            end
            begin
              dma2mem[21][26].run()  ;
            end

            begin
              gen[21][27].run()  ;
            end
            begin
              drv[21][27].run()  ;
            end
            begin
              dma2mem[21][27].run()  ;
            end

            begin
              gen[21][28].run()  ;
            end
            begin
              drv[21][28].run()  ;
            end
            begin
              dma2mem[21][28].run()  ;
            end

            begin
              gen[21][29].run()  ;
            end
            begin
              drv[21][29].run()  ;
            end
            begin
              dma2mem[21][29].run()  ;
            end

            begin
              gen[21][30].run()  ;
            end
            begin
              drv[21][30].run()  ;
            end
            begin
              dma2mem[21][30].run()  ;
            end

            begin
              gen[21][31].run()  ;
            end
            begin
              drv[21][31].run()  ;
            end
            begin
              dma2mem[21][31].run()  ;
            end

            begin
              gen[22][0].run()  ;
            end
            begin
              drv[22][0].run()  ;
            end
            begin
              dma2mem[22][0].run()  ;
            end

            begin
              gen[22][1].run()  ;
            end
            begin
              drv[22][1].run()  ;
            end
            begin
              dma2mem[22][1].run()  ;
            end

            begin
              gen[22][2].run()  ;
            end
            begin
              drv[22][2].run()  ;
            end
            begin
              dma2mem[22][2].run()  ;
            end

            begin
              gen[22][3].run()  ;
            end
            begin
              drv[22][3].run()  ;
            end
            begin
              dma2mem[22][3].run()  ;
            end

            begin
              gen[22][4].run()  ;
            end
            begin
              drv[22][4].run()  ;
            end
            begin
              dma2mem[22][4].run()  ;
            end

            begin
              gen[22][5].run()  ;
            end
            begin
              drv[22][5].run()  ;
            end
            begin
              dma2mem[22][5].run()  ;
            end

            begin
              gen[22][6].run()  ;
            end
            begin
              drv[22][6].run()  ;
            end
            begin
              dma2mem[22][6].run()  ;
            end

            begin
              gen[22][7].run()  ;
            end
            begin
              drv[22][7].run()  ;
            end
            begin
              dma2mem[22][7].run()  ;
            end

            begin
              gen[22][8].run()  ;
            end
            begin
              drv[22][8].run()  ;
            end
            begin
              dma2mem[22][8].run()  ;
            end

            begin
              gen[22][9].run()  ;
            end
            begin
              drv[22][9].run()  ;
            end
            begin
              dma2mem[22][9].run()  ;
            end

            begin
              gen[22][10].run()  ;
            end
            begin
              drv[22][10].run()  ;
            end
            begin
              dma2mem[22][10].run()  ;
            end

            begin
              gen[22][11].run()  ;
            end
            begin
              drv[22][11].run()  ;
            end
            begin
              dma2mem[22][11].run()  ;
            end

            begin
              gen[22][12].run()  ;
            end
            begin
              drv[22][12].run()  ;
            end
            begin
              dma2mem[22][12].run()  ;
            end

            begin
              gen[22][13].run()  ;
            end
            begin
              drv[22][13].run()  ;
            end
            begin
              dma2mem[22][13].run()  ;
            end

            begin
              gen[22][14].run()  ;
            end
            begin
              drv[22][14].run()  ;
            end
            begin
              dma2mem[22][14].run()  ;
            end

            begin
              gen[22][15].run()  ;
            end
            begin
              drv[22][15].run()  ;
            end
            begin
              dma2mem[22][15].run()  ;
            end

            begin
              gen[22][16].run()  ;
            end
            begin
              drv[22][16].run()  ;
            end
            begin
              dma2mem[22][16].run()  ;
            end

            begin
              gen[22][17].run()  ;
            end
            begin
              drv[22][17].run()  ;
            end
            begin
              dma2mem[22][17].run()  ;
            end

            begin
              gen[22][18].run()  ;
            end
            begin
              drv[22][18].run()  ;
            end
            begin
              dma2mem[22][18].run()  ;
            end

            begin
              gen[22][19].run()  ;
            end
            begin
              drv[22][19].run()  ;
            end
            begin
              dma2mem[22][19].run()  ;
            end

            begin
              gen[22][20].run()  ;
            end
            begin
              drv[22][20].run()  ;
            end
            begin
              dma2mem[22][20].run()  ;
            end

            begin
              gen[22][21].run()  ;
            end
            begin
              drv[22][21].run()  ;
            end
            begin
              dma2mem[22][21].run()  ;
            end

            begin
              gen[22][22].run()  ;
            end
            begin
              drv[22][22].run()  ;
            end
            begin
              dma2mem[22][22].run()  ;
            end

            begin
              gen[22][23].run()  ;
            end
            begin
              drv[22][23].run()  ;
            end
            begin
              dma2mem[22][23].run()  ;
            end

            begin
              gen[22][24].run()  ;
            end
            begin
              drv[22][24].run()  ;
            end
            begin
              dma2mem[22][24].run()  ;
            end

            begin
              gen[22][25].run()  ;
            end
            begin
              drv[22][25].run()  ;
            end
            begin
              dma2mem[22][25].run()  ;
            end

            begin
              gen[22][26].run()  ;
            end
            begin
              drv[22][26].run()  ;
            end
            begin
              dma2mem[22][26].run()  ;
            end

            begin
              gen[22][27].run()  ;
            end
            begin
              drv[22][27].run()  ;
            end
            begin
              dma2mem[22][27].run()  ;
            end

            begin
              gen[22][28].run()  ;
            end
            begin
              drv[22][28].run()  ;
            end
            begin
              dma2mem[22][28].run()  ;
            end

            begin
              gen[22][29].run()  ;
            end
            begin
              drv[22][29].run()  ;
            end
            begin
              dma2mem[22][29].run()  ;
            end

            begin
              gen[22][30].run()  ;
            end
            begin
              drv[22][30].run()  ;
            end
            begin
              dma2mem[22][30].run()  ;
            end

            begin
              gen[22][31].run()  ;
            end
            begin
              drv[22][31].run()  ;
            end
            begin
              dma2mem[22][31].run()  ;
            end

            begin
              gen[23][0].run()  ;
            end
            begin
              drv[23][0].run()  ;
            end
            begin
              dma2mem[23][0].run()  ;
            end

            begin
              gen[23][1].run()  ;
            end
            begin
              drv[23][1].run()  ;
            end
            begin
              dma2mem[23][1].run()  ;
            end

            begin
              gen[23][2].run()  ;
            end
            begin
              drv[23][2].run()  ;
            end
            begin
              dma2mem[23][2].run()  ;
            end

            begin
              gen[23][3].run()  ;
            end
            begin
              drv[23][3].run()  ;
            end
            begin
              dma2mem[23][3].run()  ;
            end

            begin
              gen[23][4].run()  ;
            end
            begin
              drv[23][4].run()  ;
            end
            begin
              dma2mem[23][4].run()  ;
            end

            begin
              gen[23][5].run()  ;
            end
            begin
              drv[23][5].run()  ;
            end
            begin
              dma2mem[23][5].run()  ;
            end

            begin
              gen[23][6].run()  ;
            end
            begin
              drv[23][6].run()  ;
            end
            begin
              dma2mem[23][6].run()  ;
            end

            begin
              gen[23][7].run()  ;
            end
            begin
              drv[23][7].run()  ;
            end
            begin
              dma2mem[23][7].run()  ;
            end

            begin
              gen[23][8].run()  ;
            end
            begin
              drv[23][8].run()  ;
            end
            begin
              dma2mem[23][8].run()  ;
            end

            begin
              gen[23][9].run()  ;
            end
            begin
              drv[23][9].run()  ;
            end
            begin
              dma2mem[23][9].run()  ;
            end

            begin
              gen[23][10].run()  ;
            end
            begin
              drv[23][10].run()  ;
            end
            begin
              dma2mem[23][10].run()  ;
            end

            begin
              gen[23][11].run()  ;
            end
            begin
              drv[23][11].run()  ;
            end
            begin
              dma2mem[23][11].run()  ;
            end

            begin
              gen[23][12].run()  ;
            end
            begin
              drv[23][12].run()  ;
            end
            begin
              dma2mem[23][12].run()  ;
            end

            begin
              gen[23][13].run()  ;
            end
            begin
              drv[23][13].run()  ;
            end
            begin
              dma2mem[23][13].run()  ;
            end

            begin
              gen[23][14].run()  ;
            end
            begin
              drv[23][14].run()  ;
            end
            begin
              dma2mem[23][14].run()  ;
            end

            begin
              gen[23][15].run()  ;
            end
            begin
              drv[23][15].run()  ;
            end
            begin
              dma2mem[23][15].run()  ;
            end

            begin
              gen[23][16].run()  ;
            end
            begin
              drv[23][16].run()  ;
            end
            begin
              dma2mem[23][16].run()  ;
            end

            begin
              gen[23][17].run()  ;
            end
            begin
              drv[23][17].run()  ;
            end
            begin
              dma2mem[23][17].run()  ;
            end

            begin
              gen[23][18].run()  ;
            end
            begin
              drv[23][18].run()  ;
            end
            begin
              dma2mem[23][18].run()  ;
            end

            begin
              gen[23][19].run()  ;
            end
            begin
              drv[23][19].run()  ;
            end
            begin
              dma2mem[23][19].run()  ;
            end

            begin
              gen[23][20].run()  ;
            end
            begin
              drv[23][20].run()  ;
            end
            begin
              dma2mem[23][20].run()  ;
            end

            begin
              gen[23][21].run()  ;
            end
            begin
              drv[23][21].run()  ;
            end
            begin
              dma2mem[23][21].run()  ;
            end

            begin
              gen[23][22].run()  ;
            end
            begin
              drv[23][22].run()  ;
            end
            begin
              dma2mem[23][22].run()  ;
            end

            begin
              gen[23][23].run()  ;
            end
            begin
              drv[23][23].run()  ;
            end
            begin
              dma2mem[23][23].run()  ;
            end

            begin
              gen[23][24].run()  ;
            end
            begin
              drv[23][24].run()  ;
            end
            begin
              dma2mem[23][24].run()  ;
            end

            begin
              gen[23][25].run()  ;
            end
            begin
              drv[23][25].run()  ;
            end
            begin
              dma2mem[23][25].run()  ;
            end

            begin
              gen[23][26].run()  ;
            end
            begin
              drv[23][26].run()  ;
            end
            begin
              dma2mem[23][26].run()  ;
            end

            begin
              gen[23][27].run()  ;
            end
            begin
              drv[23][27].run()  ;
            end
            begin
              dma2mem[23][27].run()  ;
            end

            begin
              gen[23][28].run()  ;
            end
            begin
              drv[23][28].run()  ;
            end
            begin
              dma2mem[23][28].run()  ;
            end

            begin
              gen[23][29].run()  ;
            end
            begin
              drv[23][29].run()  ;
            end
            begin
              dma2mem[23][29].run()  ;
            end

            begin
              gen[23][30].run()  ;
            end
            begin
              drv[23][30].run()  ;
            end
            begin
              dma2mem[23][30].run()  ;
            end

            begin
              gen[23][31].run()  ;
            end
            begin
              drv[23][31].run()  ;
            end
            begin
              dma2mem[23][31].run()  ;
            end

            begin
              gen[24][0].run()  ;
            end
            begin
              drv[24][0].run()  ;
            end
            begin
              dma2mem[24][0].run()  ;
            end

            begin
              gen[24][1].run()  ;
            end
            begin
              drv[24][1].run()  ;
            end
            begin
              dma2mem[24][1].run()  ;
            end

            begin
              gen[24][2].run()  ;
            end
            begin
              drv[24][2].run()  ;
            end
            begin
              dma2mem[24][2].run()  ;
            end

            begin
              gen[24][3].run()  ;
            end
            begin
              drv[24][3].run()  ;
            end
            begin
              dma2mem[24][3].run()  ;
            end

            begin
              gen[24][4].run()  ;
            end
            begin
              drv[24][4].run()  ;
            end
            begin
              dma2mem[24][4].run()  ;
            end

            begin
              gen[24][5].run()  ;
            end
            begin
              drv[24][5].run()  ;
            end
            begin
              dma2mem[24][5].run()  ;
            end

            begin
              gen[24][6].run()  ;
            end
            begin
              drv[24][6].run()  ;
            end
            begin
              dma2mem[24][6].run()  ;
            end

            begin
              gen[24][7].run()  ;
            end
            begin
              drv[24][7].run()  ;
            end
            begin
              dma2mem[24][7].run()  ;
            end

            begin
              gen[24][8].run()  ;
            end
            begin
              drv[24][8].run()  ;
            end
            begin
              dma2mem[24][8].run()  ;
            end

            begin
              gen[24][9].run()  ;
            end
            begin
              drv[24][9].run()  ;
            end
            begin
              dma2mem[24][9].run()  ;
            end

            begin
              gen[24][10].run()  ;
            end
            begin
              drv[24][10].run()  ;
            end
            begin
              dma2mem[24][10].run()  ;
            end

            begin
              gen[24][11].run()  ;
            end
            begin
              drv[24][11].run()  ;
            end
            begin
              dma2mem[24][11].run()  ;
            end

            begin
              gen[24][12].run()  ;
            end
            begin
              drv[24][12].run()  ;
            end
            begin
              dma2mem[24][12].run()  ;
            end

            begin
              gen[24][13].run()  ;
            end
            begin
              drv[24][13].run()  ;
            end
            begin
              dma2mem[24][13].run()  ;
            end

            begin
              gen[24][14].run()  ;
            end
            begin
              drv[24][14].run()  ;
            end
            begin
              dma2mem[24][14].run()  ;
            end

            begin
              gen[24][15].run()  ;
            end
            begin
              drv[24][15].run()  ;
            end
            begin
              dma2mem[24][15].run()  ;
            end

            begin
              gen[24][16].run()  ;
            end
            begin
              drv[24][16].run()  ;
            end
            begin
              dma2mem[24][16].run()  ;
            end

            begin
              gen[24][17].run()  ;
            end
            begin
              drv[24][17].run()  ;
            end
            begin
              dma2mem[24][17].run()  ;
            end

            begin
              gen[24][18].run()  ;
            end
            begin
              drv[24][18].run()  ;
            end
            begin
              dma2mem[24][18].run()  ;
            end

            begin
              gen[24][19].run()  ;
            end
            begin
              drv[24][19].run()  ;
            end
            begin
              dma2mem[24][19].run()  ;
            end

            begin
              gen[24][20].run()  ;
            end
            begin
              drv[24][20].run()  ;
            end
            begin
              dma2mem[24][20].run()  ;
            end

            begin
              gen[24][21].run()  ;
            end
            begin
              drv[24][21].run()  ;
            end
            begin
              dma2mem[24][21].run()  ;
            end

            begin
              gen[24][22].run()  ;
            end
            begin
              drv[24][22].run()  ;
            end
            begin
              dma2mem[24][22].run()  ;
            end

            begin
              gen[24][23].run()  ;
            end
            begin
              drv[24][23].run()  ;
            end
            begin
              dma2mem[24][23].run()  ;
            end

            begin
              gen[24][24].run()  ;
            end
            begin
              drv[24][24].run()  ;
            end
            begin
              dma2mem[24][24].run()  ;
            end

            begin
              gen[24][25].run()  ;
            end
            begin
              drv[24][25].run()  ;
            end
            begin
              dma2mem[24][25].run()  ;
            end

            begin
              gen[24][26].run()  ;
            end
            begin
              drv[24][26].run()  ;
            end
            begin
              dma2mem[24][26].run()  ;
            end

            begin
              gen[24][27].run()  ;
            end
            begin
              drv[24][27].run()  ;
            end
            begin
              dma2mem[24][27].run()  ;
            end

            begin
              gen[24][28].run()  ;
            end
            begin
              drv[24][28].run()  ;
            end
            begin
              dma2mem[24][28].run()  ;
            end

            begin
              gen[24][29].run()  ;
            end
            begin
              drv[24][29].run()  ;
            end
            begin
              dma2mem[24][29].run()  ;
            end

            begin
              gen[24][30].run()  ;
            end
            begin
              drv[24][30].run()  ;
            end
            begin
              dma2mem[24][30].run()  ;
            end

            begin
              gen[24][31].run()  ;
            end
            begin
              drv[24][31].run()  ;
            end
            begin
              dma2mem[24][31].run()  ;
            end

            begin
              gen[25][0].run()  ;
            end
            begin
              drv[25][0].run()  ;
            end
            begin
              dma2mem[25][0].run()  ;
            end

            begin
              gen[25][1].run()  ;
            end
            begin
              drv[25][1].run()  ;
            end
            begin
              dma2mem[25][1].run()  ;
            end

            begin
              gen[25][2].run()  ;
            end
            begin
              drv[25][2].run()  ;
            end
            begin
              dma2mem[25][2].run()  ;
            end

            begin
              gen[25][3].run()  ;
            end
            begin
              drv[25][3].run()  ;
            end
            begin
              dma2mem[25][3].run()  ;
            end

            begin
              gen[25][4].run()  ;
            end
            begin
              drv[25][4].run()  ;
            end
            begin
              dma2mem[25][4].run()  ;
            end

            begin
              gen[25][5].run()  ;
            end
            begin
              drv[25][5].run()  ;
            end
            begin
              dma2mem[25][5].run()  ;
            end

            begin
              gen[25][6].run()  ;
            end
            begin
              drv[25][6].run()  ;
            end
            begin
              dma2mem[25][6].run()  ;
            end

            begin
              gen[25][7].run()  ;
            end
            begin
              drv[25][7].run()  ;
            end
            begin
              dma2mem[25][7].run()  ;
            end

            begin
              gen[25][8].run()  ;
            end
            begin
              drv[25][8].run()  ;
            end
            begin
              dma2mem[25][8].run()  ;
            end

            begin
              gen[25][9].run()  ;
            end
            begin
              drv[25][9].run()  ;
            end
            begin
              dma2mem[25][9].run()  ;
            end

            begin
              gen[25][10].run()  ;
            end
            begin
              drv[25][10].run()  ;
            end
            begin
              dma2mem[25][10].run()  ;
            end

            begin
              gen[25][11].run()  ;
            end
            begin
              drv[25][11].run()  ;
            end
            begin
              dma2mem[25][11].run()  ;
            end

            begin
              gen[25][12].run()  ;
            end
            begin
              drv[25][12].run()  ;
            end
            begin
              dma2mem[25][12].run()  ;
            end

            begin
              gen[25][13].run()  ;
            end
            begin
              drv[25][13].run()  ;
            end
            begin
              dma2mem[25][13].run()  ;
            end

            begin
              gen[25][14].run()  ;
            end
            begin
              drv[25][14].run()  ;
            end
            begin
              dma2mem[25][14].run()  ;
            end

            begin
              gen[25][15].run()  ;
            end
            begin
              drv[25][15].run()  ;
            end
            begin
              dma2mem[25][15].run()  ;
            end

            begin
              gen[25][16].run()  ;
            end
            begin
              drv[25][16].run()  ;
            end
            begin
              dma2mem[25][16].run()  ;
            end

            begin
              gen[25][17].run()  ;
            end
            begin
              drv[25][17].run()  ;
            end
            begin
              dma2mem[25][17].run()  ;
            end

            begin
              gen[25][18].run()  ;
            end
            begin
              drv[25][18].run()  ;
            end
            begin
              dma2mem[25][18].run()  ;
            end

            begin
              gen[25][19].run()  ;
            end
            begin
              drv[25][19].run()  ;
            end
            begin
              dma2mem[25][19].run()  ;
            end

            begin
              gen[25][20].run()  ;
            end
            begin
              drv[25][20].run()  ;
            end
            begin
              dma2mem[25][20].run()  ;
            end

            begin
              gen[25][21].run()  ;
            end
            begin
              drv[25][21].run()  ;
            end
            begin
              dma2mem[25][21].run()  ;
            end

            begin
              gen[25][22].run()  ;
            end
            begin
              drv[25][22].run()  ;
            end
            begin
              dma2mem[25][22].run()  ;
            end

            begin
              gen[25][23].run()  ;
            end
            begin
              drv[25][23].run()  ;
            end
            begin
              dma2mem[25][23].run()  ;
            end

            begin
              gen[25][24].run()  ;
            end
            begin
              drv[25][24].run()  ;
            end
            begin
              dma2mem[25][24].run()  ;
            end

            begin
              gen[25][25].run()  ;
            end
            begin
              drv[25][25].run()  ;
            end
            begin
              dma2mem[25][25].run()  ;
            end

            begin
              gen[25][26].run()  ;
            end
            begin
              drv[25][26].run()  ;
            end
            begin
              dma2mem[25][26].run()  ;
            end

            begin
              gen[25][27].run()  ;
            end
            begin
              drv[25][27].run()  ;
            end
            begin
              dma2mem[25][27].run()  ;
            end

            begin
              gen[25][28].run()  ;
            end
            begin
              drv[25][28].run()  ;
            end
            begin
              dma2mem[25][28].run()  ;
            end

            begin
              gen[25][29].run()  ;
            end
            begin
              drv[25][29].run()  ;
            end
            begin
              dma2mem[25][29].run()  ;
            end

            begin
              gen[25][30].run()  ;
            end
            begin
              drv[25][30].run()  ;
            end
            begin
              dma2mem[25][30].run()  ;
            end

            begin
              gen[25][31].run()  ;
            end
            begin
              drv[25][31].run()  ;
            end
            begin
              dma2mem[25][31].run()  ;
            end

            begin
              gen[26][0].run()  ;
            end
            begin
              drv[26][0].run()  ;
            end
            begin
              dma2mem[26][0].run()  ;
            end

            begin
              gen[26][1].run()  ;
            end
            begin
              drv[26][1].run()  ;
            end
            begin
              dma2mem[26][1].run()  ;
            end

            begin
              gen[26][2].run()  ;
            end
            begin
              drv[26][2].run()  ;
            end
            begin
              dma2mem[26][2].run()  ;
            end

            begin
              gen[26][3].run()  ;
            end
            begin
              drv[26][3].run()  ;
            end
            begin
              dma2mem[26][3].run()  ;
            end

            begin
              gen[26][4].run()  ;
            end
            begin
              drv[26][4].run()  ;
            end
            begin
              dma2mem[26][4].run()  ;
            end

            begin
              gen[26][5].run()  ;
            end
            begin
              drv[26][5].run()  ;
            end
            begin
              dma2mem[26][5].run()  ;
            end

            begin
              gen[26][6].run()  ;
            end
            begin
              drv[26][6].run()  ;
            end
            begin
              dma2mem[26][6].run()  ;
            end

            begin
              gen[26][7].run()  ;
            end
            begin
              drv[26][7].run()  ;
            end
            begin
              dma2mem[26][7].run()  ;
            end

            begin
              gen[26][8].run()  ;
            end
            begin
              drv[26][8].run()  ;
            end
            begin
              dma2mem[26][8].run()  ;
            end

            begin
              gen[26][9].run()  ;
            end
            begin
              drv[26][9].run()  ;
            end
            begin
              dma2mem[26][9].run()  ;
            end

            begin
              gen[26][10].run()  ;
            end
            begin
              drv[26][10].run()  ;
            end
            begin
              dma2mem[26][10].run()  ;
            end

            begin
              gen[26][11].run()  ;
            end
            begin
              drv[26][11].run()  ;
            end
            begin
              dma2mem[26][11].run()  ;
            end

            begin
              gen[26][12].run()  ;
            end
            begin
              drv[26][12].run()  ;
            end
            begin
              dma2mem[26][12].run()  ;
            end

            begin
              gen[26][13].run()  ;
            end
            begin
              drv[26][13].run()  ;
            end
            begin
              dma2mem[26][13].run()  ;
            end

            begin
              gen[26][14].run()  ;
            end
            begin
              drv[26][14].run()  ;
            end
            begin
              dma2mem[26][14].run()  ;
            end

            begin
              gen[26][15].run()  ;
            end
            begin
              drv[26][15].run()  ;
            end
            begin
              dma2mem[26][15].run()  ;
            end

            begin
              gen[26][16].run()  ;
            end
            begin
              drv[26][16].run()  ;
            end
            begin
              dma2mem[26][16].run()  ;
            end

            begin
              gen[26][17].run()  ;
            end
            begin
              drv[26][17].run()  ;
            end
            begin
              dma2mem[26][17].run()  ;
            end

            begin
              gen[26][18].run()  ;
            end
            begin
              drv[26][18].run()  ;
            end
            begin
              dma2mem[26][18].run()  ;
            end

            begin
              gen[26][19].run()  ;
            end
            begin
              drv[26][19].run()  ;
            end
            begin
              dma2mem[26][19].run()  ;
            end

            begin
              gen[26][20].run()  ;
            end
            begin
              drv[26][20].run()  ;
            end
            begin
              dma2mem[26][20].run()  ;
            end

            begin
              gen[26][21].run()  ;
            end
            begin
              drv[26][21].run()  ;
            end
            begin
              dma2mem[26][21].run()  ;
            end

            begin
              gen[26][22].run()  ;
            end
            begin
              drv[26][22].run()  ;
            end
            begin
              dma2mem[26][22].run()  ;
            end

            begin
              gen[26][23].run()  ;
            end
            begin
              drv[26][23].run()  ;
            end
            begin
              dma2mem[26][23].run()  ;
            end

            begin
              gen[26][24].run()  ;
            end
            begin
              drv[26][24].run()  ;
            end
            begin
              dma2mem[26][24].run()  ;
            end

            begin
              gen[26][25].run()  ;
            end
            begin
              drv[26][25].run()  ;
            end
            begin
              dma2mem[26][25].run()  ;
            end

            begin
              gen[26][26].run()  ;
            end
            begin
              drv[26][26].run()  ;
            end
            begin
              dma2mem[26][26].run()  ;
            end

            begin
              gen[26][27].run()  ;
            end
            begin
              drv[26][27].run()  ;
            end
            begin
              dma2mem[26][27].run()  ;
            end

            begin
              gen[26][28].run()  ;
            end
            begin
              drv[26][28].run()  ;
            end
            begin
              dma2mem[26][28].run()  ;
            end

            begin
              gen[26][29].run()  ;
            end
            begin
              drv[26][29].run()  ;
            end
            begin
              dma2mem[26][29].run()  ;
            end

            begin
              gen[26][30].run()  ;
            end
            begin
              drv[26][30].run()  ;
            end
            begin
              dma2mem[26][30].run()  ;
            end

            begin
              gen[26][31].run()  ;
            end
            begin
              drv[26][31].run()  ;
            end
            begin
              dma2mem[26][31].run()  ;
            end

            begin
              gen[27][0].run()  ;
            end
            begin
              drv[27][0].run()  ;
            end
            begin
              dma2mem[27][0].run()  ;
            end

            begin
              gen[27][1].run()  ;
            end
            begin
              drv[27][1].run()  ;
            end
            begin
              dma2mem[27][1].run()  ;
            end

            begin
              gen[27][2].run()  ;
            end
            begin
              drv[27][2].run()  ;
            end
            begin
              dma2mem[27][2].run()  ;
            end

            begin
              gen[27][3].run()  ;
            end
            begin
              drv[27][3].run()  ;
            end
            begin
              dma2mem[27][3].run()  ;
            end

            begin
              gen[27][4].run()  ;
            end
            begin
              drv[27][4].run()  ;
            end
            begin
              dma2mem[27][4].run()  ;
            end

            begin
              gen[27][5].run()  ;
            end
            begin
              drv[27][5].run()  ;
            end
            begin
              dma2mem[27][5].run()  ;
            end

            begin
              gen[27][6].run()  ;
            end
            begin
              drv[27][6].run()  ;
            end
            begin
              dma2mem[27][6].run()  ;
            end

            begin
              gen[27][7].run()  ;
            end
            begin
              drv[27][7].run()  ;
            end
            begin
              dma2mem[27][7].run()  ;
            end

            begin
              gen[27][8].run()  ;
            end
            begin
              drv[27][8].run()  ;
            end
            begin
              dma2mem[27][8].run()  ;
            end

            begin
              gen[27][9].run()  ;
            end
            begin
              drv[27][9].run()  ;
            end
            begin
              dma2mem[27][9].run()  ;
            end

            begin
              gen[27][10].run()  ;
            end
            begin
              drv[27][10].run()  ;
            end
            begin
              dma2mem[27][10].run()  ;
            end

            begin
              gen[27][11].run()  ;
            end
            begin
              drv[27][11].run()  ;
            end
            begin
              dma2mem[27][11].run()  ;
            end

            begin
              gen[27][12].run()  ;
            end
            begin
              drv[27][12].run()  ;
            end
            begin
              dma2mem[27][12].run()  ;
            end

            begin
              gen[27][13].run()  ;
            end
            begin
              drv[27][13].run()  ;
            end
            begin
              dma2mem[27][13].run()  ;
            end

            begin
              gen[27][14].run()  ;
            end
            begin
              drv[27][14].run()  ;
            end
            begin
              dma2mem[27][14].run()  ;
            end

            begin
              gen[27][15].run()  ;
            end
            begin
              drv[27][15].run()  ;
            end
            begin
              dma2mem[27][15].run()  ;
            end

            begin
              gen[27][16].run()  ;
            end
            begin
              drv[27][16].run()  ;
            end
            begin
              dma2mem[27][16].run()  ;
            end

            begin
              gen[27][17].run()  ;
            end
            begin
              drv[27][17].run()  ;
            end
            begin
              dma2mem[27][17].run()  ;
            end

            begin
              gen[27][18].run()  ;
            end
            begin
              drv[27][18].run()  ;
            end
            begin
              dma2mem[27][18].run()  ;
            end

            begin
              gen[27][19].run()  ;
            end
            begin
              drv[27][19].run()  ;
            end
            begin
              dma2mem[27][19].run()  ;
            end

            begin
              gen[27][20].run()  ;
            end
            begin
              drv[27][20].run()  ;
            end
            begin
              dma2mem[27][20].run()  ;
            end

            begin
              gen[27][21].run()  ;
            end
            begin
              drv[27][21].run()  ;
            end
            begin
              dma2mem[27][21].run()  ;
            end

            begin
              gen[27][22].run()  ;
            end
            begin
              drv[27][22].run()  ;
            end
            begin
              dma2mem[27][22].run()  ;
            end

            begin
              gen[27][23].run()  ;
            end
            begin
              drv[27][23].run()  ;
            end
            begin
              dma2mem[27][23].run()  ;
            end

            begin
              gen[27][24].run()  ;
            end
            begin
              drv[27][24].run()  ;
            end
            begin
              dma2mem[27][24].run()  ;
            end

            begin
              gen[27][25].run()  ;
            end
            begin
              drv[27][25].run()  ;
            end
            begin
              dma2mem[27][25].run()  ;
            end

            begin
              gen[27][26].run()  ;
            end
            begin
              drv[27][26].run()  ;
            end
            begin
              dma2mem[27][26].run()  ;
            end

            begin
              gen[27][27].run()  ;
            end
            begin
              drv[27][27].run()  ;
            end
            begin
              dma2mem[27][27].run()  ;
            end

            begin
              gen[27][28].run()  ;
            end
            begin
              drv[27][28].run()  ;
            end
            begin
              dma2mem[27][28].run()  ;
            end

            begin
              gen[27][29].run()  ;
            end
            begin
              drv[27][29].run()  ;
            end
            begin
              dma2mem[27][29].run()  ;
            end

            begin
              gen[27][30].run()  ;
            end
            begin
              drv[27][30].run()  ;
            end
            begin
              dma2mem[27][30].run()  ;
            end

            begin
              gen[27][31].run()  ;
            end
            begin
              drv[27][31].run()  ;
            end
            begin
              dma2mem[27][31].run()  ;
            end

            begin
              gen[28][0].run()  ;
            end
            begin
              drv[28][0].run()  ;
            end
            begin
              dma2mem[28][0].run()  ;
            end

            begin
              gen[28][1].run()  ;
            end
            begin
              drv[28][1].run()  ;
            end
            begin
              dma2mem[28][1].run()  ;
            end

            begin
              gen[28][2].run()  ;
            end
            begin
              drv[28][2].run()  ;
            end
            begin
              dma2mem[28][2].run()  ;
            end

            begin
              gen[28][3].run()  ;
            end
            begin
              drv[28][3].run()  ;
            end
            begin
              dma2mem[28][3].run()  ;
            end

            begin
              gen[28][4].run()  ;
            end
            begin
              drv[28][4].run()  ;
            end
            begin
              dma2mem[28][4].run()  ;
            end

            begin
              gen[28][5].run()  ;
            end
            begin
              drv[28][5].run()  ;
            end
            begin
              dma2mem[28][5].run()  ;
            end

            begin
              gen[28][6].run()  ;
            end
            begin
              drv[28][6].run()  ;
            end
            begin
              dma2mem[28][6].run()  ;
            end

            begin
              gen[28][7].run()  ;
            end
            begin
              drv[28][7].run()  ;
            end
            begin
              dma2mem[28][7].run()  ;
            end

            begin
              gen[28][8].run()  ;
            end
            begin
              drv[28][8].run()  ;
            end
            begin
              dma2mem[28][8].run()  ;
            end

            begin
              gen[28][9].run()  ;
            end
            begin
              drv[28][9].run()  ;
            end
            begin
              dma2mem[28][9].run()  ;
            end

            begin
              gen[28][10].run()  ;
            end
            begin
              drv[28][10].run()  ;
            end
            begin
              dma2mem[28][10].run()  ;
            end

            begin
              gen[28][11].run()  ;
            end
            begin
              drv[28][11].run()  ;
            end
            begin
              dma2mem[28][11].run()  ;
            end

            begin
              gen[28][12].run()  ;
            end
            begin
              drv[28][12].run()  ;
            end
            begin
              dma2mem[28][12].run()  ;
            end

            begin
              gen[28][13].run()  ;
            end
            begin
              drv[28][13].run()  ;
            end
            begin
              dma2mem[28][13].run()  ;
            end

            begin
              gen[28][14].run()  ;
            end
            begin
              drv[28][14].run()  ;
            end
            begin
              dma2mem[28][14].run()  ;
            end

            begin
              gen[28][15].run()  ;
            end
            begin
              drv[28][15].run()  ;
            end
            begin
              dma2mem[28][15].run()  ;
            end

            begin
              gen[28][16].run()  ;
            end
            begin
              drv[28][16].run()  ;
            end
            begin
              dma2mem[28][16].run()  ;
            end

            begin
              gen[28][17].run()  ;
            end
            begin
              drv[28][17].run()  ;
            end
            begin
              dma2mem[28][17].run()  ;
            end

            begin
              gen[28][18].run()  ;
            end
            begin
              drv[28][18].run()  ;
            end
            begin
              dma2mem[28][18].run()  ;
            end

            begin
              gen[28][19].run()  ;
            end
            begin
              drv[28][19].run()  ;
            end
            begin
              dma2mem[28][19].run()  ;
            end

            begin
              gen[28][20].run()  ;
            end
            begin
              drv[28][20].run()  ;
            end
            begin
              dma2mem[28][20].run()  ;
            end

            begin
              gen[28][21].run()  ;
            end
            begin
              drv[28][21].run()  ;
            end
            begin
              dma2mem[28][21].run()  ;
            end

            begin
              gen[28][22].run()  ;
            end
            begin
              drv[28][22].run()  ;
            end
            begin
              dma2mem[28][22].run()  ;
            end

            begin
              gen[28][23].run()  ;
            end
            begin
              drv[28][23].run()  ;
            end
            begin
              dma2mem[28][23].run()  ;
            end

            begin
              gen[28][24].run()  ;
            end
            begin
              drv[28][24].run()  ;
            end
            begin
              dma2mem[28][24].run()  ;
            end

            begin
              gen[28][25].run()  ;
            end
            begin
              drv[28][25].run()  ;
            end
            begin
              dma2mem[28][25].run()  ;
            end

            begin
              gen[28][26].run()  ;
            end
            begin
              drv[28][26].run()  ;
            end
            begin
              dma2mem[28][26].run()  ;
            end

            begin
              gen[28][27].run()  ;
            end
            begin
              drv[28][27].run()  ;
            end
            begin
              dma2mem[28][27].run()  ;
            end

            begin
              gen[28][28].run()  ;
            end
            begin
              drv[28][28].run()  ;
            end
            begin
              dma2mem[28][28].run()  ;
            end

            begin
              gen[28][29].run()  ;
            end
            begin
              drv[28][29].run()  ;
            end
            begin
              dma2mem[28][29].run()  ;
            end

            begin
              gen[28][30].run()  ;
            end
            begin
              drv[28][30].run()  ;
            end
            begin
              dma2mem[28][30].run()  ;
            end

            begin
              gen[28][31].run()  ;
            end
            begin
              drv[28][31].run()  ;
            end
            begin
              dma2mem[28][31].run()  ;
            end

            begin
              gen[29][0].run()  ;
            end
            begin
              drv[29][0].run()  ;
            end
            begin
              dma2mem[29][0].run()  ;
            end

            begin
              gen[29][1].run()  ;
            end
            begin
              drv[29][1].run()  ;
            end
            begin
              dma2mem[29][1].run()  ;
            end

            begin
              gen[29][2].run()  ;
            end
            begin
              drv[29][2].run()  ;
            end
            begin
              dma2mem[29][2].run()  ;
            end

            begin
              gen[29][3].run()  ;
            end
            begin
              drv[29][3].run()  ;
            end
            begin
              dma2mem[29][3].run()  ;
            end

            begin
              gen[29][4].run()  ;
            end
            begin
              drv[29][4].run()  ;
            end
            begin
              dma2mem[29][4].run()  ;
            end

            begin
              gen[29][5].run()  ;
            end
            begin
              drv[29][5].run()  ;
            end
            begin
              dma2mem[29][5].run()  ;
            end

            begin
              gen[29][6].run()  ;
            end
            begin
              drv[29][6].run()  ;
            end
            begin
              dma2mem[29][6].run()  ;
            end

            begin
              gen[29][7].run()  ;
            end
            begin
              drv[29][7].run()  ;
            end
            begin
              dma2mem[29][7].run()  ;
            end

            begin
              gen[29][8].run()  ;
            end
            begin
              drv[29][8].run()  ;
            end
            begin
              dma2mem[29][8].run()  ;
            end

            begin
              gen[29][9].run()  ;
            end
            begin
              drv[29][9].run()  ;
            end
            begin
              dma2mem[29][9].run()  ;
            end

            begin
              gen[29][10].run()  ;
            end
            begin
              drv[29][10].run()  ;
            end
            begin
              dma2mem[29][10].run()  ;
            end

            begin
              gen[29][11].run()  ;
            end
            begin
              drv[29][11].run()  ;
            end
            begin
              dma2mem[29][11].run()  ;
            end

            begin
              gen[29][12].run()  ;
            end
            begin
              drv[29][12].run()  ;
            end
            begin
              dma2mem[29][12].run()  ;
            end

            begin
              gen[29][13].run()  ;
            end
            begin
              drv[29][13].run()  ;
            end
            begin
              dma2mem[29][13].run()  ;
            end

            begin
              gen[29][14].run()  ;
            end
            begin
              drv[29][14].run()  ;
            end
            begin
              dma2mem[29][14].run()  ;
            end

            begin
              gen[29][15].run()  ;
            end
            begin
              drv[29][15].run()  ;
            end
            begin
              dma2mem[29][15].run()  ;
            end

            begin
              gen[29][16].run()  ;
            end
            begin
              drv[29][16].run()  ;
            end
            begin
              dma2mem[29][16].run()  ;
            end

            begin
              gen[29][17].run()  ;
            end
            begin
              drv[29][17].run()  ;
            end
            begin
              dma2mem[29][17].run()  ;
            end

            begin
              gen[29][18].run()  ;
            end
            begin
              drv[29][18].run()  ;
            end
            begin
              dma2mem[29][18].run()  ;
            end

            begin
              gen[29][19].run()  ;
            end
            begin
              drv[29][19].run()  ;
            end
            begin
              dma2mem[29][19].run()  ;
            end

            begin
              gen[29][20].run()  ;
            end
            begin
              drv[29][20].run()  ;
            end
            begin
              dma2mem[29][20].run()  ;
            end

            begin
              gen[29][21].run()  ;
            end
            begin
              drv[29][21].run()  ;
            end
            begin
              dma2mem[29][21].run()  ;
            end

            begin
              gen[29][22].run()  ;
            end
            begin
              drv[29][22].run()  ;
            end
            begin
              dma2mem[29][22].run()  ;
            end

            begin
              gen[29][23].run()  ;
            end
            begin
              drv[29][23].run()  ;
            end
            begin
              dma2mem[29][23].run()  ;
            end

            begin
              gen[29][24].run()  ;
            end
            begin
              drv[29][24].run()  ;
            end
            begin
              dma2mem[29][24].run()  ;
            end

            begin
              gen[29][25].run()  ;
            end
            begin
              drv[29][25].run()  ;
            end
            begin
              dma2mem[29][25].run()  ;
            end

            begin
              gen[29][26].run()  ;
            end
            begin
              drv[29][26].run()  ;
            end
            begin
              dma2mem[29][26].run()  ;
            end

            begin
              gen[29][27].run()  ;
            end
            begin
              drv[29][27].run()  ;
            end
            begin
              dma2mem[29][27].run()  ;
            end

            begin
              gen[29][28].run()  ;
            end
            begin
              drv[29][28].run()  ;
            end
            begin
              dma2mem[29][28].run()  ;
            end

            begin
              gen[29][29].run()  ;
            end
            begin
              drv[29][29].run()  ;
            end
            begin
              dma2mem[29][29].run()  ;
            end

            begin
              gen[29][30].run()  ;
            end
            begin
              drv[29][30].run()  ;
            end
            begin
              dma2mem[29][30].run()  ;
            end

            begin
              gen[29][31].run()  ;
            end
            begin
              drv[29][31].run()  ;
            end
            begin
              dma2mem[29][31].run()  ;
            end

            begin
              gen[30][0].run()  ;
            end
            begin
              drv[30][0].run()  ;
            end
            begin
              dma2mem[30][0].run()  ;
            end

            begin
              gen[30][1].run()  ;
            end
            begin
              drv[30][1].run()  ;
            end
            begin
              dma2mem[30][1].run()  ;
            end

            begin
              gen[30][2].run()  ;
            end
            begin
              drv[30][2].run()  ;
            end
            begin
              dma2mem[30][2].run()  ;
            end

            begin
              gen[30][3].run()  ;
            end
            begin
              drv[30][3].run()  ;
            end
            begin
              dma2mem[30][3].run()  ;
            end

            begin
              gen[30][4].run()  ;
            end
            begin
              drv[30][4].run()  ;
            end
            begin
              dma2mem[30][4].run()  ;
            end

            begin
              gen[30][5].run()  ;
            end
            begin
              drv[30][5].run()  ;
            end
            begin
              dma2mem[30][5].run()  ;
            end

            begin
              gen[30][6].run()  ;
            end
            begin
              drv[30][6].run()  ;
            end
            begin
              dma2mem[30][6].run()  ;
            end

            begin
              gen[30][7].run()  ;
            end
            begin
              drv[30][7].run()  ;
            end
            begin
              dma2mem[30][7].run()  ;
            end

            begin
              gen[30][8].run()  ;
            end
            begin
              drv[30][8].run()  ;
            end
            begin
              dma2mem[30][8].run()  ;
            end

            begin
              gen[30][9].run()  ;
            end
            begin
              drv[30][9].run()  ;
            end
            begin
              dma2mem[30][9].run()  ;
            end

            begin
              gen[30][10].run()  ;
            end
            begin
              drv[30][10].run()  ;
            end
            begin
              dma2mem[30][10].run()  ;
            end

            begin
              gen[30][11].run()  ;
            end
            begin
              drv[30][11].run()  ;
            end
            begin
              dma2mem[30][11].run()  ;
            end

            begin
              gen[30][12].run()  ;
            end
            begin
              drv[30][12].run()  ;
            end
            begin
              dma2mem[30][12].run()  ;
            end

            begin
              gen[30][13].run()  ;
            end
            begin
              drv[30][13].run()  ;
            end
            begin
              dma2mem[30][13].run()  ;
            end

            begin
              gen[30][14].run()  ;
            end
            begin
              drv[30][14].run()  ;
            end
            begin
              dma2mem[30][14].run()  ;
            end

            begin
              gen[30][15].run()  ;
            end
            begin
              drv[30][15].run()  ;
            end
            begin
              dma2mem[30][15].run()  ;
            end

            begin
              gen[30][16].run()  ;
            end
            begin
              drv[30][16].run()  ;
            end
            begin
              dma2mem[30][16].run()  ;
            end

            begin
              gen[30][17].run()  ;
            end
            begin
              drv[30][17].run()  ;
            end
            begin
              dma2mem[30][17].run()  ;
            end

            begin
              gen[30][18].run()  ;
            end
            begin
              drv[30][18].run()  ;
            end
            begin
              dma2mem[30][18].run()  ;
            end

            begin
              gen[30][19].run()  ;
            end
            begin
              drv[30][19].run()  ;
            end
            begin
              dma2mem[30][19].run()  ;
            end

            begin
              gen[30][20].run()  ;
            end
            begin
              drv[30][20].run()  ;
            end
            begin
              dma2mem[30][20].run()  ;
            end

            begin
              gen[30][21].run()  ;
            end
            begin
              drv[30][21].run()  ;
            end
            begin
              dma2mem[30][21].run()  ;
            end

            begin
              gen[30][22].run()  ;
            end
            begin
              drv[30][22].run()  ;
            end
            begin
              dma2mem[30][22].run()  ;
            end

            begin
              gen[30][23].run()  ;
            end
            begin
              drv[30][23].run()  ;
            end
            begin
              dma2mem[30][23].run()  ;
            end

            begin
              gen[30][24].run()  ;
            end
            begin
              drv[30][24].run()  ;
            end
            begin
              dma2mem[30][24].run()  ;
            end

            begin
              gen[30][25].run()  ;
            end
            begin
              drv[30][25].run()  ;
            end
            begin
              dma2mem[30][25].run()  ;
            end

            begin
              gen[30][26].run()  ;
            end
            begin
              drv[30][26].run()  ;
            end
            begin
              dma2mem[30][26].run()  ;
            end

            begin
              gen[30][27].run()  ;
            end
            begin
              drv[30][27].run()  ;
            end
            begin
              dma2mem[30][27].run()  ;
            end

            begin
              gen[30][28].run()  ;
            end
            begin
              drv[30][28].run()  ;
            end
            begin
              dma2mem[30][28].run()  ;
            end

            begin
              gen[30][29].run()  ;
            end
            begin
              drv[30][29].run()  ;
            end
            begin
              dma2mem[30][29].run()  ;
            end

            begin
              gen[30][30].run()  ;
            end
            begin
              drv[30][30].run()  ;
            end
            begin
              dma2mem[30][30].run()  ;
            end

            begin
              gen[30][31].run()  ;
            end
            begin
              drv[30][31].run()  ;
            end
            begin
              dma2mem[30][31].run()  ;
            end

            begin
              gen[31][0].run()  ;
            end
            begin
              drv[31][0].run()  ;
            end
            begin
              dma2mem[31][0].run()  ;
            end

            begin
              gen[31][1].run()  ;
            end
            begin
              drv[31][1].run()  ;
            end
            begin
              dma2mem[31][1].run()  ;
            end

            begin
              gen[31][2].run()  ;
            end
            begin
              drv[31][2].run()  ;
            end
            begin
              dma2mem[31][2].run()  ;
            end

            begin
              gen[31][3].run()  ;
            end
            begin
              drv[31][3].run()  ;
            end
            begin
              dma2mem[31][3].run()  ;
            end

            begin
              gen[31][4].run()  ;
            end
            begin
              drv[31][4].run()  ;
            end
            begin
              dma2mem[31][4].run()  ;
            end

            begin
              gen[31][5].run()  ;
            end
            begin
              drv[31][5].run()  ;
            end
            begin
              dma2mem[31][5].run()  ;
            end

            begin
              gen[31][6].run()  ;
            end
            begin
              drv[31][6].run()  ;
            end
            begin
              dma2mem[31][6].run()  ;
            end

            begin
              gen[31][7].run()  ;
            end
            begin
              drv[31][7].run()  ;
            end
            begin
              dma2mem[31][7].run()  ;
            end

            begin
              gen[31][8].run()  ;
            end
            begin
              drv[31][8].run()  ;
            end
            begin
              dma2mem[31][8].run()  ;
            end

            begin
              gen[31][9].run()  ;
            end
            begin
              drv[31][9].run()  ;
            end
            begin
              dma2mem[31][9].run()  ;
            end

            begin
              gen[31][10].run()  ;
            end
            begin
              drv[31][10].run()  ;
            end
            begin
              dma2mem[31][10].run()  ;
            end

            begin
              gen[31][11].run()  ;
            end
            begin
              drv[31][11].run()  ;
            end
            begin
              dma2mem[31][11].run()  ;
            end

            begin
              gen[31][12].run()  ;
            end
            begin
              drv[31][12].run()  ;
            end
            begin
              dma2mem[31][12].run()  ;
            end

            begin
              gen[31][13].run()  ;
            end
            begin
              drv[31][13].run()  ;
            end
            begin
              dma2mem[31][13].run()  ;
            end

            begin
              gen[31][14].run()  ;
            end
            begin
              drv[31][14].run()  ;
            end
            begin
              dma2mem[31][14].run()  ;
            end

            begin
              gen[31][15].run()  ;
            end
            begin
              drv[31][15].run()  ;
            end
            begin
              dma2mem[31][15].run()  ;
            end

            begin
              gen[31][16].run()  ;
            end
            begin
              drv[31][16].run()  ;
            end
            begin
              dma2mem[31][16].run()  ;
            end

            begin
              gen[31][17].run()  ;
            end
            begin
              drv[31][17].run()  ;
            end
            begin
              dma2mem[31][17].run()  ;
            end

            begin
              gen[31][18].run()  ;
            end
            begin
              drv[31][18].run()  ;
            end
            begin
              dma2mem[31][18].run()  ;
            end

            begin
              gen[31][19].run()  ;
            end
            begin
              drv[31][19].run()  ;
            end
            begin
              dma2mem[31][19].run()  ;
            end

            begin
              gen[31][20].run()  ;
            end
            begin
              drv[31][20].run()  ;
            end
            begin
              dma2mem[31][20].run()  ;
            end

            begin
              gen[31][21].run()  ;
            end
            begin
              drv[31][21].run()  ;
            end
            begin
              dma2mem[31][21].run()  ;
            end

            begin
              gen[31][22].run()  ;
            end
            begin
              drv[31][22].run()  ;
            end
            begin
              dma2mem[31][22].run()  ;
            end

            begin
              gen[31][23].run()  ;
            end
            begin
              drv[31][23].run()  ;
            end
            begin
              dma2mem[31][23].run()  ;
            end

            begin
              gen[31][24].run()  ;
            end
            begin
              drv[31][24].run()  ;
            end
            begin
              dma2mem[31][24].run()  ;
            end

            begin
              gen[31][25].run()  ;
            end
            begin
              drv[31][25].run()  ;
            end
            begin
              dma2mem[31][25].run()  ;
            end

            begin
              gen[31][26].run()  ;
            end
            begin
              drv[31][26].run()  ;
            end
            begin
              dma2mem[31][26].run()  ;
            end

            begin
              gen[31][27].run()  ;
            end
            begin
              drv[31][27].run()  ;
            end
            begin
              dma2mem[31][27].run()  ;
            end

            begin
              gen[31][28].run()  ;
            end
            begin
              drv[31][28].run()  ;
            end
            begin
              dma2mem[31][28].run()  ;
            end

            begin
              gen[31][29].run()  ;
            end
            begin
              drv[31][29].run()  ;
            end
            begin
              dma2mem[31][29].run()  ;
            end

            begin
              gen[31][30].run()  ;
            end
            begin
              drv[31][30].run()  ;
            end
            begin
              dma2mem[31][30].run()  ;
            end

            begin
              gen[31][31].run()  ;
            end
            begin
              drv[31][31].run()  ;
            end
            begin
              dma2mem[31][31].run()  ;
            end

            begin
              gen[32][0].run()  ;
            end
            begin
              drv[32][0].run()  ;
            end
            begin
              dma2mem[32][0].run()  ;
            end

            begin
              gen[32][1].run()  ;
            end
            begin
              drv[32][1].run()  ;
            end
            begin
              dma2mem[32][1].run()  ;
            end

            begin
              gen[32][2].run()  ;
            end
            begin
              drv[32][2].run()  ;
            end
            begin
              dma2mem[32][2].run()  ;
            end

            begin
              gen[32][3].run()  ;
            end
            begin
              drv[32][3].run()  ;
            end
            begin
              dma2mem[32][3].run()  ;
            end

            begin
              gen[32][4].run()  ;
            end
            begin
              drv[32][4].run()  ;
            end
            begin
              dma2mem[32][4].run()  ;
            end

            begin
              gen[32][5].run()  ;
            end
            begin
              drv[32][5].run()  ;
            end
            begin
              dma2mem[32][5].run()  ;
            end

            begin
              gen[32][6].run()  ;
            end
            begin
              drv[32][6].run()  ;
            end
            begin
              dma2mem[32][6].run()  ;
            end

            begin
              gen[32][7].run()  ;
            end
            begin
              drv[32][7].run()  ;
            end
            begin
              dma2mem[32][7].run()  ;
            end

            begin
              gen[32][8].run()  ;
            end
            begin
              drv[32][8].run()  ;
            end
            begin
              dma2mem[32][8].run()  ;
            end

            begin
              gen[32][9].run()  ;
            end
            begin
              drv[32][9].run()  ;
            end
            begin
              dma2mem[32][9].run()  ;
            end

            begin
              gen[32][10].run()  ;
            end
            begin
              drv[32][10].run()  ;
            end
            begin
              dma2mem[32][10].run()  ;
            end

            begin
              gen[32][11].run()  ;
            end
            begin
              drv[32][11].run()  ;
            end
            begin
              dma2mem[32][11].run()  ;
            end

            begin
              gen[32][12].run()  ;
            end
            begin
              drv[32][12].run()  ;
            end
            begin
              dma2mem[32][12].run()  ;
            end

            begin
              gen[32][13].run()  ;
            end
            begin
              drv[32][13].run()  ;
            end
            begin
              dma2mem[32][13].run()  ;
            end

            begin
              gen[32][14].run()  ;
            end
            begin
              drv[32][14].run()  ;
            end
            begin
              dma2mem[32][14].run()  ;
            end

            begin
              gen[32][15].run()  ;
            end
            begin
              drv[32][15].run()  ;
            end
            begin
              dma2mem[32][15].run()  ;
            end

            begin
              gen[32][16].run()  ;
            end
            begin
              drv[32][16].run()  ;
            end
            begin
              dma2mem[32][16].run()  ;
            end

            begin
              gen[32][17].run()  ;
            end
            begin
              drv[32][17].run()  ;
            end
            begin
              dma2mem[32][17].run()  ;
            end

            begin
              gen[32][18].run()  ;
            end
            begin
              drv[32][18].run()  ;
            end
            begin
              dma2mem[32][18].run()  ;
            end

            begin
              gen[32][19].run()  ;
            end
            begin
              drv[32][19].run()  ;
            end
            begin
              dma2mem[32][19].run()  ;
            end

            begin
              gen[32][20].run()  ;
            end
            begin
              drv[32][20].run()  ;
            end
            begin
              dma2mem[32][20].run()  ;
            end

            begin
              gen[32][21].run()  ;
            end
            begin
              drv[32][21].run()  ;
            end
            begin
              dma2mem[32][21].run()  ;
            end

            begin
              gen[32][22].run()  ;
            end
            begin
              drv[32][22].run()  ;
            end
            begin
              dma2mem[32][22].run()  ;
            end

            begin
              gen[32][23].run()  ;
            end
            begin
              drv[32][23].run()  ;
            end
            begin
              dma2mem[32][23].run()  ;
            end

            begin
              gen[32][24].run()  ;
            end
            begin
              drv[32][24].run()  ;
            end
            begin
              dma2mem[32][24].run()  ;
            end

            begin
              gen[32][25].run()  ;
            end
            begin
              drv[32][25].run()  ;
            end
            begin
              dma2mem[32][25].run()  ;
            end

            begin
              gen[32][26].run()  ;
            end
            begin
              drv[32][26].run()  ;
            end
            begin
              dma2mem[32][26].run()  ;
            end

            begin
              gen[32][27].run()  ;
            end
            begin
              drv[32][27].run()  ;
            end
            begin
              dma2mem[32][27].run()  ;
            end

            begin
              gen[32][28].run()  ;
            end
            begin
              drv[32][28].run()  ;
            end
            begin
              dma2mem[32][28].run()  ;
            end

            begin
              gen[32][29].run()  ;
            end
            begin
              drv[32][29].run()  ;
            end
            begin
              dma2mem[32][29].run()  ;
            end

            begin
              gen[32][30].run()  ;
            end
            begin
              drv[32][30].run()  ;
            end
            begin
              dma2mem[32][30].run()  ;
            end

            begin
              gen[32][31].run()  ;
            end
            begin
              drv[32][31].run()  ;
            end
            begin
              dma2mem[32][31].run()  ;
            end

            begin
              gen[33][0].run()  ;
            end
            begin
              drv[33][0].run()  ;
            end
            begin
              dma2mem[33][0].run()  ;
            end

            begin
              gen[33][1].run()  ;
            end
            begin
              drv[33][1].run()  ;
            end
            begin
              dma2mem[33][1].run()  ;
            end

            begin
              gen[33][2].run()  ;
            end
            begin
              drv[33][2].run()  ;
            end
            begin
              dma2mem[33][2].run()  ;
            end

            begin
              gen[33][3].run()  ;
            end
            begin
              drv[33][3].run()  ;
            end
            begin
              dma2mem[33][3].run()  ;
            end

            begin
              gen[33][4].run()  ;
            end
            begin
              drv[33][4].run()  ;
            end
            begin
              dma2mem[33][4].run()  ;
            end

            begin
              gen[33][5].run()  ;
            end
            begin
              drv[33][5].run()  ;
            end
            begin
              dma2mem[33][5].run()  ;
            end

            begin
              gen[33][6].run()  ;
            end
            begin
              drv[33][6].run()  ;
            end
            begin
              dma2mem[33][6].run()  ;
            end

            begin
              gen[33][7].run()  ;
            end
            begin
              drv[33][7].run()  ;
            end
            begin
              dma2mem[33][7].run()  ;
            end

            begin
              gen[33][8].run()  ;
            end
            begin
              drv[33][8].run()  ;
            end
            begin
              dma2mem[33][8].run()  ;
            end

            begin
              gen[33][9].run()  ;
            end
            begin
              drv[33][9].run()  ;
            end
            begin
              dma2mem[33][9].run()  ;
            end

            begin
              gen[33][10].run()  ;
            end
            begin
              drv[33][10].run()  ;
            end
            begin
              dma2mem[33][10].run()  ;
            end

            begin
              gen[33][11].run()  ;
            end
            begin
              drv[33][11].run()  ;
            end
            begin
              dma2mem[33][11].run()  ;
            end

            begin
              gen[33][12].run()  ;
            end
            begin
              drv[33][12].run()  ;
            end
            begin
              dma2mem[33][12].run()  ;
            end

            begin
              gen[33][13].run()  ;
            end
            begin
              drv[33][13].run()  ;
            end
            begin
              dma2mem[33][13].run()  ;
            end

            begin
              gen[33][14].run()  ;
            end
            begin
              drv[33][14].run()  ;
            end
            begin
              dma2mem[33][14].run()  ;
            end

            begin
              gen[33][15].run()  ;
            end
            begin
              drv[33][15].run()  ;
            end
            begin
              dma2mem[33][15].run()  ;
            end

            begin
              gen[33][16].run()  ;
            end
            begin
              drv[33][16].run()  ;
            end
            begin
              dma2mem[33][16].run()  ;
            end

            begin
              gen[33][17].run()  ;
            end
            begin
              drv[33][17].run()  ;
            end
            begin
              dma2mem[33][17].run()  ;
            end

            begin
              gen[33][18].run()  ;
            end
            begin
              drv[33][18].run()  ;
            end
            begin
              dma2mem[33][18].run()  ;
            end

            begin
              gen[33][19].run()  ;
            end
            begin
              drv[33][19].run()  ;
            end
            begin
              dma2mem[33][19].run()  ;
            end

            begin
              gen[33][20].run()  ;
            end
            begin
              drv[33][20].run()  ;
            end
            begin
              dma2mem[33][20].run()  ;
            end

            begin
              gen[33][21].run()  ;
            end
            begin
              drv[33][21].run()  ;
            end
            begin
              dma2mem[33][21].run()  ;
            end

            begin
              gen[33][22].run()  ;
            end
            begin
              drv[33][22].run()  ;
            end
            begin
              dma2mem[33][22].run()  ;
            end

            begin
              gen[33][23].run()  ;
            end
            begin
              drv[33][23].run()  ;
            end
            begin
              dma2mem[33][23].run()  ;
            end

            begin
              gen[33][24].run()  ;
            end
            begin
              drv[33][24].run()  ;
            end
            begin
              dma2mem[33][24].run()  ;
            end

            begin
              gen[33][25].run()  ;
            end
            begin
              drv[33][25].run()  ;
            end
            begin
              dma2mem[33][25].run()  ;
            end

            begin
              gen[33][26].run()  ;
            end
            begin
              drv[33][26].run()  ;
            end
            begin
              dma2mem[33][26].run()  ;
            end

            begin
              gen[33][27].run()  ;
            end
            begin
              drv[33][27].run()  ;
            end
            begin
              dma2mem[33][27].run()  ;
            end

            begin
              gen[33][28].run()  ;
            end
            begin
              drv[33][28].run()  ;
            end
            begin
              dma2mem[33][28].run()  ;
            end

            begin
              gen[33][29].run()  ;
            end
            begin
              drv[33][29].run()  ;
            end
            begin
              dma2mem[33][29].run()  ;
            end

            begin
              gen[33][30].run()  ;
            end
            begin
              drv[33][30].run()  ;
            end
            begin
              dma2mem[33][30].run()  ;
            end

            begin
              gen[33][31].run()  ;
            end
            begin
              drv[33][31].run()  ;
            end
            begin
              dma2mem[33][31].run()  ;
            end

            begin
              gen[34][0].run()  ;
            end
            begin
              drv[34][0].run()  ;
            end
            begin
              dma2mem[34][0].run()  ;
            end

            begin
              gen[34][1].run()  ;
            end
            begin
              drv[34][1].run()  ;
            end
            begin
              dma2mem[34][1].run()  ;
            end

            begin
              gen[34][2].run()  ;
            end
            begin
              drv[34][2].run()  ;
            end
            begin
              dma2mem[34][2].run()  ;
            end

            begin
              gen[34][3].run()  ;
            end
            begin
              drv[34][3].run()  ;
            end
            begin
              dma2mem[34][3].run()  ;
            end

            begin
              gen[34][4].run()  ;
            end
            begin
              drv[34][4].run()  ;
            end
            begin
              dma2mem[34][4].run()  ;
            end

            begin
              gen[34][5].run()  ;
            end
            begin
              drv[34][5].run()  ;
            end
            begin
              dma2mem[34][5].run()  ;
            end

            begin
              gen[34][6].run()  ;
            end
            begin
              drv[34][6].run()  ;
            end
            begin
              dma2mem[34][6].run()  ;
            end

            begin
              gen[34][7].run()  ;
            end
            begin
              drv[34][7].run()  ;
            end
            begin
              dma2mem[34][7].run()  ;
            end

            begin
              gen[34][8].run()  ;
            end
            begin
              drv[34][8].run()  ;
            end
            begin
              dma2mem[34][8].run()  ;
            end

            begin
              gen[34][9].run()  ;
            end
            begin
              drv[34][9].run()  ;
            end
            begin
              dma2mem[34][9].run()  ;
            end

            begin
              gen[34][10].run()  ;
            end
            begin
              drv[34][10].run()  ;
            end
            begin
              dma2mem[34][10].run()  ;
            end

            begin
              gen[34][11].run()  ;
            end
            begin
              drv[34][11].run()  ;
            end
            begin
              dma2mem[34][11].run()  ;
            end

            begin
              gen[34][12].run()  ;
            end
            begin
              drv[34][12].run()  ;
            end
            begin
              dma2mem[34][12].run()  ;
            end

            begin
              gen[34][13].run()  ;
            end
            begin
              drv[34][13].run()  ;
            end
            begin
              dma2mem[34][13].run()  ;
            end

            begin
              gen[34][14].run()  ;
            end
            begin
              drv[34][14].run()  ;
            end
            begin
              dma2mem[34][14].run()  ;
            end

            begin
              gen[34][15].run()  ;
            end
            begin
              drv[34][15].run()  ;
            end
            begin
              dma2mem[34][15].run()  ;
            end

            begin
              gen[34][16].run()  ;
            end
            begin
              drv[34][16].run()  ;
            end
            begin
              dma2mem[34][16].run()  ;
            end

            begin
              gen[34][17].run()  ;
            end
            begin
              drv[34][17].run()  ;
            end
            begin
              dma2mem[34][17].run()  ;
            end

            begin
              gen[34][18].run()  ;
            end
            begin
              drv[34][18].run()  ;
            end
            begin
              dma2mem[34][18].run()  ;
            end

            begin
              gen[34][19].run()  ;
            end
            begin
              drv[34][19].run()  ;
            end
            begin
              dma2mem[34][19].run()  ;
            end

            begin
              gen[34][20].run()  ;
            end
            begin
              drv[34][20].run()  ;
            end
            begin
              dma2mem[34][20].run()  ;
            end

            begin
              gen[34][21].run()  ;
            end
            begin
              drv[34][21].run()  ;
            end
            begin
              dma2mem[34][21].run()  ;
            end

            begin
              gen[34][22].run()  ;
            end
            begin
              drv[34][22].run()  ;
            end
            begin
              dma2mem[34][22].run()  ;
            end

            begin
              gen[34][23].run()  ;
            end
            begin
              drv[34][23].run()  ;
            end
            begin
              dma2mem[34][23].run()  ;
            end

            begin
              gen[34][24].run()  ;
            end
            begin
              drv[34][24].run()  ;
            end
            begin
              dma2mem[34][24].run()  ;
            end

            begin
              gen[34][25].run()  ;
            end
            begin
              drv[34][25].run()  ;
            end
            begin
              dma2mem[34][25].run()  ;
            end

            begin
              gen[34][26].run()  ;
            end
            begin
              drv[34][26].run()  ;
            end
            begin
              dma2mem[34][26].run()  ;
            end

            begin
              gen[34][27].run()  ;
            end
            begin
              drv[34][27].run()  ;
            end
            begin
              dma2mem[34][27].run()  ;
            end

            begin
              gen[34][28].run()  ;
            end
            begin
              drv[34][28].run()  ;
            end
            begin
              dma2mem[34][28].run()  ;
            end

            begin
              gen[34][29].run()  ;
            end
            begin
              drv[34][29].run()  ;
            end
            begin
              dma2mem[34][29].run()  ;
            end

            begin
              gen[34][30].run()  ;
            end
            begin
              drv[34][30].run()  ;
            end
            begin
              dma2mem[34][30].run()  ;
            end

            begin
              gen[34][31].run()  ;
            end
            begin
              drv[34][31].run()  ;
            end
            begin
              dma2mem[34][31].run()  ;
            end

            begin
              gen[35][0].run()  ;
            end
            begin
              drv[35][0].run()  ;
            end
            begin
              dma2mem[35][0].run()  ;
            end

            begin
              gen[35][1].run()  ;
            end
            begin
              drv[35][1].run()  ;
            end
            begin
              dma2mem[35][1].run()  ;
            end

            begin
              gen[35][2].run()  ;
            end
            begin
              drv[35][2].run()  ;
            end
            begin
              dma2mem[35][2].run()  ;
            end

            begin
              gen[35][3].run()  ;
            end
            begin
              drv[35][3].run()  ;
            end
            begin
              dma2mem[35][3].run()  ;
            end

            begin
              gen[35][4].run()  ;
            end
            begin
              drv[35][4].run()  ;
            end
            begin
              dma2mem[35][4].run()  ;
            end

            begin
              gen[35][5].run()  ;
            end
            begin
              drv[35][5].run()  ;
            end
            begin
              dma2mem[35][5].run()  ;
            end

            begin
              gen[35][6].run()  ;
            end
            begin
              drv[35][6].run()  ;
            end
            begin
              dma2mem[35][6].run()  ;
            end

            begin
              gen[35][7].run()  ;
            end
            begin
              drv[35][7].run()  ;
            end
            begin
              dma2mem[35][7].run()  ;
            end

            begin
              gen[35][8].run()  ;
            end
            begin
              drv[35][8].run()  ;
            end
            begin
              dma2mem[35][8].run()  ;
            end

            begin
              gen[35][9].run()  ;
            end
            begin
              drv[35][9].run()  ;
            end
            begin
              dma2mem[35][9].run()  ;
            end

            begin
              gen[35][10].run()  ;
            end
            begin
              drv[35][10].run()  ;
            end
            begin
              dma2mem[35][10].run()  ;
            end

            begin
              gen[35][11].run()  ;
            end
            begin
              drv[35][11].run()  ;
            end
            begin
              dma2mem[35][11].run()  ;
            end

            begin
              gen[35][12].run()  ;
            end
            begin
              drv[35][12].run()  ;
            end
            begin
              dma2mem[35][12].run()  ;
            end

            begin
              gen[35][13].run()  ;
            end
            begin
              drv[35][13].run()  ;
            end
            begin
              dma2mem[35][13].run()  ;
            end

            begin
              gen[35][14].run()  ;
            end
            begin
              drv[35][14].run()  ;
            end
            begin
              dma2mem[35][14].run()  ;
            end

            begin
              gen[35][15].run()  ;
            end
            begin
              drv[35][15].run()  ;
            end
            begin
              dma2mem[35][15].run()  ;
            end

            begin
              gen[35][16].run()  ;
            end
            begin
              drv[35][16].run()  ;
            end
            begin
              dma2mem[35][16].run()  ;
            end

            begin
              gen[35][17].run()  ;
            end
            begin
              drv[35][17].run()  ;
            end
            begin
              dma2mem[35][17].run()  ;
            end

            begin
              gen[35][18].run()  ;
            end
            begin
              drv[35][18].run()  ;
            end
            begin
              dma2mem[35][18].run()  ;
            end

            begin
              gen[35][19].run()  ;
            end
            begin
              drv[35][19].run()  ;
            end
            begin
              dma2mem[35][19].run()  ;
            end

            begin
              gen[35][20].run()  ;
            end
            begin
              drv[35][20].run()  ;
            end
            begin
              dma2mem[35][20].run()  ;
            end

            begin
              gen[35][21].run()  ;
            end
            begin
              drv[35][21].run()  ;
            end
            begin
              dma2mem[35][21].run()  ;
            end

            begin
              gen[35][22].run()  ;
            end
            begin
              drv[35][22].run()  ;
            end
            begin
              dma2mem[35][22].run()  ;
            end

            begin
              gen[35][23].run()  ;
            end
            begin
              drv[35][23].run()  ;
            end
            begin
              dma2mem[35][23].run()  ;
            end

            begin
              gen[35][24].run()  ;
            end
            begin
              drv[35][24].run()  ;
            end
            begin
              dma2mem[35][24].run()  ;
            end

            begin
              gen[35][25].run()  ;
            end
            begin
              drv[35][25].run()  ;
            end
            begin
              dma2mem[35][25].run()  ;
            end

            begin
              gen[35][26].run()  ;
            end
            begin
              drv[35][26].run()  ;
            end
            begin
              dma2mem[35][26].run()  ;
            end

            begin
              gen[35][27].run()  ;
            end
            begin
              drv[35][27].run()  ;
            end
            begin
              dma2mem[35][27].run()  ;
            end

            begin
              gen[35][28].run()  ;
            end
            begin
              drv[35][28].run()  ;
            end
            begin
              dma2mem[35][28].run()  ;
            end

            begin
              gen[35][29].run()  ;
            end
            begin
              drv[35][29].run()  ;
            end
            begin
              dma2mem[35][29].run()  ;
            end

            begin
              gen[35][30].run()  ;
            end
            begin
              drv[35][30].run()  ;
            end
            begin
              dma2mem[35][30].run()  ;
            end

            begin
              gen[35][31].run()  ;
            end
            begin
              drv[35][31].run()  ;
            end
            begin
              dma2mem[35][31].run()  ;
            end

            begin
              gen[36][0].run()  ;
            end
            begin
              drv[36][0].run()  ;
            end
            begin
              dma2mem[36][0].run()  ;
            end

            begin
              gen[36][1].run()  ;
            end
            begin
              drv[36][1].run()  ;
            end
            begin
              dma2mem[36][1].run()  ;
            end

            begin
              gen[36][2].run()  ;
            end
            begin
              drv[36][2].run()  ;
            end
            begin
              dma2mem[36][2].run()  ;
            end

            begin
              gen[36][3].run()  ;
            end
            begin
              drv[36][3].run()  ;
            end
            begin
              dma2mem[36][3].run()  ;
            end

            begin
              gen[36][4].run()  ;
            end
            begin
              drv[36][4].run()  ;
            end
            begin
              dma2mem[36][4].run()  ;
            end

            begin
              gen[36][5].run()  ;
            end
            begin
              drv[36][5].run()  ;
            end
            begin
              dma2mem[36][5].run()  ;
            end

            begin
              gen[36][6].run()  ;
            end
            begin
              drv[36][6].run()  ;
            end
            begin
              dma2mem[36][6].run()  ;
            end

            begin
              gen[36][7].run()  ;
            end
            begin
              drv[36][7].run()  ;
            end
            begin
              dma2mem[36][7].run()  ;
            end

            begin
              gen[36][8].run()  ;
            end
            begin
              drv[36][8].run()  ;
            end
            begin
              dma2mem[36][8].run()  ;
            end

            begin
              gen[36][9].run()  ;
            end
            begin
              drv[36][9].run()  ;
            end
            begin
              dma2mem[36][9].run()  ;
            end

            begin
              gen[36][10].run()  ;
            end
            begin
              drv[36][10].run()  ;
            end
            begin
              dma2mem[36][10].run()  ;
            end

            begin
              gen[36][11].run()  ;
            end
            begin
              drv[36][11].run()  ;
            end
            begin
              dma2mem[36][11].run()  ;
            end

            begin
              gen[36][12].run()  ;
            end
            begin
              drv[36][12].run()  ;
            end
            begin
              dma2mem[36][12].run()  ;
            end

            begin
              gen[36][13].run()  ;
            end
            begin
              drv[36][13].run()  ;
            end
            begin
              dma2mem[36][13].run()  ;
            end

            begin
              gen[36][14].run()  ;
            end
            begin
              drv[36][14].run()  ;
            end
            begin
              dma2mem[36][14].run()  ;
            end

            begin
              gen[36][15].run()  ;
            end
            begin
              drv[36][15].run()  ;
            end
            begin
              dma2mem[36][15].run()  ;
            end

            begin
              gen[36][16].run()  ;
            end
            begin
              drv[36][16].run()  ;
            end
            begin
              dma2mem[36][16].run()  ;
            end

            begin
              gen[36][17].run()  ;
            end
            begin
              drv[36][17].run()  ;
            end
            begin
              dma2mem[36][17].run()  ;
            end

            begin
              gen[36][18].run()  ;
            end
            begin
              drv[36][18].run()  ;
            end
            begin
              dma2mem[36][18].run()  ;
            end

            begin
              gen[36][19].run()  ;
            end
            begin
              drv[36][19].run()  ;
            end
            begin
              dma2mem[36][19].run()  ;
            end

            begin
              gen[36][20].run()  ;
            end
            begin
              drv[36][20].run()  ;
            end
            begin
              dma2mem[36][20].run()  ;
            end

            begin
              gen[36][21].run()  ;
            end
            begin
              drv[36][21].run()  ;
            end
            begin
              dma2mem[36][21].run()  ;
            end

            begin
              gen[36][22].run()  ;
            end
            begin
              drv[36][22].run()  ;
            end
            begin
              dma2mem[36][22].run()  ;
            end

            begin
              gen[36][23].run()  ;
            end
            begin
              drv[36][23].run()  ;
            end
            begin
              dma2mem[36][23].run()  ;
            end

            begin
              gen[36][24].run()  ;
            end
            begin
              drv[36][24].run()  ;
            end
            begin
              dma2mem[36][24].run()  ;
            end

            begin
              gen[36][25].run()  ;
            end
            begin
              drv[36][25].run()  ;
            end
            begin
              dma2mem[36][25].run()  ;
            end

            begin
              gen[36][26].run()  ;
            end
            begin
              drv[36][26].run()  ;
            end
            begin
              dma2mem[36][26].run()  ;
            end

            begin
              gen[36][27].run()  ;
            end
            begin
              drv[36][27].run()  ;
            end
            begin
              dma2mem[36][27].run()  ;
            end

            begin
              gen[36][28].run()  ;
            end
            begin
              drv[36][28].run()  ;
            end
            begin
              dma2mem[36][28].run()  ;
            end

            begin
              gen[36][29].run()  ;
            end
            begin
              drv[36][29].run()  ;
            end
            begin
              dma2mem[36][29].run()  ;
            end

            begin
              gen[36][30].run()  ;
            end
            begin
              drv[36][30].run()  ;
            end
            begin
              dma2mem[36][30].run()  ;
            end

            begin
              gen[36][31].run()  ;
            end
            begin
              drv[36][31].run()  ;
            end
            begin
              dma2mem[36][31].run()  ;
            end

            begin
              gen[37][0].run()  ;
            end
            begin
              drv[37][0].run()  ;
            end
            begin
              dma2mem[37][0].run()  ;
            end

            begin
              gen[37][1].run()  ;
            end
            begin
              drv[37][1].run()  ;
            end
            begin
              dma2mem[37][1].run()  ;
            end

            begin
              gen[37][2].run()  ;
            end
            begin
              drv[37][2].run()  ;
            end
            begin
              dma2mem[37][2].run()  ;
            end

            begin
              gen[37][3].run()  ;
            end
            begin
              drv[37][3].run()  ;
            end
            begin
              dma2mem[37][3].run()  ;
            end

            begin
              gen[37][4].run()  ;
            end
            begin
              drv[37][4].run()  ;
            end
            begin
              dma2mem[37][4].run()  ;
            end

            begin
              gen[37][5].run()  ;
            end
            begin
              drv[37][5].run()  ;
            end
            begin
              dma2mem[37][5].run()  ;
            end

            begin
              gen[37][6].run()  ;
            end
            begin
              drv[37][6].run()  ;
            end
            begin
              dma2mem[37][6].run()  ;
            end

            begin
              gen[37][7].run()  ;
            end
            begin
              drv[37][7].run()  ;
            end
            begin
              dma2mem[37][7].run()  ;
            end

            begin
              gen[37][8].run()  ;
            end
            begin
              drv[37][8].run()  ;
            end
            begin
              dma2mem[37][8].run()  ;
            end

            begin
              gen[37][9].run()  ;
            end
            begin
              drv[37][9].run()  ;
            end
            begin
              dma2mem[37][9].run()  ;
            end

            begin
              gen[37][10].run()  ;
            end
            begin
              drv[37][10].run()  ;
            end
            begin
              dma2mem[37][10].run()  ;
            end

            begin
              gen[37][11].run()  ;
            end
            begin
              drv[37][11].run()  ;
            end
            begin
              dma2mem[37][11].run()  ;
            end

            begin
              gen[37][12].run()  ;
            end
            begin
              drv[37][12].run()  ;
            end
            begin
              dma2mem[37][12].run()  ;
            end

            begin
              gen[37][13].run()  ;
            end
            begin
              drv[37][13].run()  ;
            end
            begin
              dma2mem[37][13].run()  ;
            end

            begin
              gen[37][14].run()  ;
            end
            begin
              drv[37][14].run()  ;
            end
            begin
              dma2mem[37][14].run()  ;
            end

            begin
              gen[37][15].run()  ;
            end
            begin
              drv[37][15].run()  ;
            end
            begin
              dma2mem[37][15].run()  ;
            end

            begin
              gen[37][16].run()  ;
            end
            begin
              drv[37][16].run()  ;
            end
            begin
              dma2mem[37][16].run()  ;
            end

            begin
              gen[37][17].run()  ;
            end
            begin
              drv[37][17].run()  ;
            end
            begin
              dma2mem[37][17].run()  ;
            end

            begin
              gen[37][18].run()  ;
            end
            begin
              drv[37][18].run()  ;
            end
            begin
              dma2mem[37][18].run()  ;
            end

            begin
              gen[37][19].run()  ;
            end
            begin
              drv[37][19].run()  ;
            end
            begin
              dma2mem[37][19].run()  ;
            end

            begin
              gen[37][20].run()  ;
            end
            begin
              drv[37][20].run()  ;
            end
            begin
              dma2mem[37][20].run()  ;
            end

            begin
              gen[37][21].run()  ;
            end
            begin
              drv[37][21].run()  ;
            end
            begin
              dma2mem[37][21].run()  ;
            end

            begin
              gen[37][22].run()  ;
            end
            begin
              drv[37][22].run()  ;
            end
            begin
              dma2mem[37][22].run()  ;
            end

            begin
              gen[37][23].run()  ;
            end
            begin
              drv[37][23].run()  ;
            end
            begin
              dma2mem[37][23].run()  ;
            end

            begin
              gen[37][24].run()  ;
            end
            begin
              drv[37][24].run()  ;
            end
            begin
              dma2mem[37][24].run()  ;
            end

            begin
              gen[37][25].run()  ;
            end
            begin
              drv[37][25].run()  ;
            end
            begin
              dma2mem[37][25].run()  ;
            end

            begin
              gen[37][26].run()  ;
            end
            begin
              drv[37][26].run()  ;
            end
            begin
              dma2mem[37][26].run()  ;
            end

            begin
              gen[37][27].run()  ;
            end
            begin
              drv[37][27].run()  ;
            end
            begin
              dma2mem[37][27].run()  ;
            end

            begin
              gen[37][28].run()  ;
            end
            begin
              drv[37][28].run()  ;
            end
            begin
              dma2mem[37][28].run()  ;
            end

            begin
              gen[37][29].run()  ;
            end
            begin
              drv[37][29].run()  ;
            end
            begin
              dma2mem[37][29].run()  ;
            end

            begin
              gen[37][30].run()  ;
            end
            begin
              drv[37][30].run()  ;
            end
            begin
              dma2mem[37][30].run()  ;
            end

            begin
              gen[37][31].run()  ;
            end
            begin
              drv[37][31].run()  ;
            end
            begin
              dma2mem[37][31].run()  ;
            end

            begin
              gen[38][0].run()  ;
            end
            begin
              drv[38][0].run()  ;
            end
            begin
              dma2mem[38][0].run()  ;
            end

            begin
              gen[38][1].run()  ;
            end
            begin
              drv[38][1].run()  ;
            end
            begin
              dma2mem[38][1].run()  ;
            end

            begin
              gen[38][2].run()  ;
            end
            begin
              drv[38][2].run()  ;
            end
            begin
              dma2mem[38][2].run()  ;
            end

            begin
              gen[38][3].run()  ;
            end
            begin
              drv[38][3].run()  ;
            end
            begin
              dma2mem[38][3].run()  ;
            end

            begin
              gen[38][4].run()  ;
            end
            begin
              drv[38][4].run()  ;
            end
            begin
              dma2mem[38][4].run()  ;
            end

            begin
              gen[38][5].run()  ;
            end
            begin
              drv[38][5].run()  ;
            end
            begin
              dma2mem[38][5].run()  ;
            end

            begin
              gen[38][6].run()  ;
            end
            begin
              drv[38][6].run()  ;
            end
            begin
              dma2mem[38][6].run()  ;
            end

            begin
              gen[38][7].run()  ;
            end
            begin
              drv[38][7].run()  ;
            end
            begin
              dma2mem[38][7].run()  ;
            end

            begin
              gen[38][8].run()  ;
            end
            begin
              drv[38][8].run()  ;
            end
            begin
              dma2mem[38][8].run()  ;
            end

            begin
              gen[38][9].run()  ;
            end
            begin
              drv[38][9].run()  ;
            end
            begin
              dma2mem[38][9].run()  ;
            end

            begin
              gen[38][10].run()  ;
            end
            begin
              drv[38][10].run()  ;
            end
            begin
              dma2mem[38][10].run()  ;
            end

            begin
              gen[38][11].run()  ;
            end
            begin
              drv[38][11].run()  ;
            end
            begin
              dma2mem[38][11].run()  ;
            end

            begin
              gen[38][12].run()  ;
            end
            begin
              drv[38][12].run()  ;
            end
            begin
              dma2mem[38][12].run()  ;
            end

            begin
              gen[38][13].run()  ;
            end
            begin
              drv[38][13].run()  ;
            end
            begin
              dma2mem[38][13].run()  ;
            end

            begin
              gen[38][14].run()  ;
            end
            begin
              drv[38][14].run()  ;
            end
            begin
              dma2mem[38][14].run()  ;
            end

            begin
              gen[38][15].run()  ;
            end
            begin
              drv[38][15].run()  ;
            end
            begin
              dma2mem[38][15].run()  ;
            end

            begin
              gen[38][16].run()  ;
            end
            begin
              drv[38][16].run()  ;
            end
            begin
              dma2mem[38][16].run()  ;
            end

            begin
              gen[38][17].run()  ;
            end
            begin
              drv[38][17].run()  ;
            end
            begin
              dma2mem[38][17].run()  ;
            end

            begin
              gen[38][18].run()  ;
            end
            begin
              drv[38][18].run()  ;
            end
            begin
              dma2mem[38][18].run()  ;
            end

            begin
              gen[38][19].run()  ;
            end
            begin
              drv[38][19].run()  ;
            end
            begin
              dma2mem[38][19].run()  ;
            end

            begin
              gen[38][20].run()  ;
            end
            begin
              drv[38][20].run()  ;
            end
            begin
              dma2mem[38][20].run()  ;
            end

            begin
              gen[38][21].run()  ;
            end
            begin
              drv[38][21].run()  ;
            end
            begin
              dma2mem[38][21].run()  ;
            end

            begin
              gen[38][22].run()  ;
            end
            begin
              drv[38][22].run()  ;
            end
            begin
              dma2mem[38][22].run()  ;
            end

            begin
              gen[38][23].run()  ;
            end
            begin
              drv[38][23].run()  ;
            end
            begin
              dma2mem[38][23].run()  ;
            end

            begin
              gen[38][24].run()  ;
            end
            begin
              drv[38][24].run()  ;
            end
            begin
              dma2mem[38][24].run()  ;
            end

            begin
              gen[38][25].run()  ;
            end
            begin
              drv[38][25].run()  ;
            end
            begin
              dma2mem[38][25].run()  ;
            end

            begin
              gen[38][26].run()  ;
            end
            begin
              drv[38][26].run()  ;
            end
            begin
              dma2mem[38][26].run()  ;
            end

            begin
              gen[38][27].run()  ;
            end
            begin
              drv[38][27].run()  ;
            end
            begin
              dma2mem[38][27].run()  ;
            end

            begin
              gen[38][28].run()  ;
            end
            begin
              drv[38][28].run()  ;
            end
            begin
              dma2mem[38][28].run()  ;
            end

            begin
              gen[38][29].run()  ;
            end
            begin
              drv[38][29].run()  ;
            end
            begin
              dma2mem[38][29].run()  ;
            end

            begin
              gen[38][30].run()  ;
            end
            begin
              drv[38][30].run()  ;
            end
            begin
              dma2mem[38][30].run()  ;
            end

            begin
              gen[38][31].run()  ;
            end
            begin
              drv[38][31].run()  ;
            end
            begin
              dma2mem[38][31].run()  ;
            end

            begin
              gen[39][0].run()  ;
            end
            begin
              drv[39][0].run()  ;
            end
            begin
              dma2mem[39][0].run()  ;
            end

            begin
              gen[39][1].run()  ;
            end
            begin
              drv[39][1].run()  ;
            end
            begin
              dma2mem[39][1].run()  ;
            end

            begin
              gen[39][2].run()  ;
            end
            begin
              drv[39][2].run()  ;
            end
            begin
              dma2mem[39][2].run()  ;
            end

            begin
              gen[39][3].run()  ;
            end
            begin
              drv[39][3].run()  ;
            end
            begin
              dma2mem[39][3].run()  ;
            end

            begin
              gen[39][4].run()  ;
            end
            begin
              drv[39][4].run()  ;
            end
            begin
              dma2mem[39][4].run()  ;
            end

            begin
              gen[39][5].run()  ;
            end
            begin
              drv[39][5].run()  ;
            end
            begin
              dma2mem[39][5].run()  ;
            end

            begin
              gen[39][6].run()  ;
            end
            begin
              drv[39][6].run()  ;
            end
            begin
              dma2mem[39][6].run()  ;
            end

            begin
              gen[39][7].run()  ;
            end
            begin
              drv[39][7].run()  ;
            end
            begin
              dma2mem[39][7].run()  ;
            end

            begin
              gen[39][8].run()  ;
            end
            begin
              drv[39][8].run()  ;
            end
            begin
              dma2mem[39][8].run()  ;
            end

            begin
              gen[39][9].run()  ;
            end
            begin
              drv[39][9].run()  ;
            end
            begin
              dma2mem[39][9].run()  ;
            end

            begin
              gen[39][10].run()  ;
            end
            begin
              drv[39][10].run()  ;
            end
            begin
              dma2mem[39][10].run()  ;
            end

            begin
              gen[39][11].run()  ;
            end
            begin
              drv[39][11].run()  ;
            end
            begin
              dma2mem[39][11].run()  ;
            end

            begin
              gen[39][12].run()  ;
            end
            begin
              drv[39][12].run()  ;
            end
            begin
              dma2mem[39][12].run()  ;
            end

            begin
              gen[39][13].run()  ;
            end
            begin
              drv[39][13].run()  ;
            end
            begin
              dma2mem[39][13].run()  ;
            end

            begin
              gen[39][14].run()  ;
            end
            begin
              drv[39][14].run()  ;
            end
            begin
              dma2mem[39][14].run()  ;
            end

            begin
              gen[39][15].run()  ;
            end
            begin
              drv[39][15].run()  ;
            end
            begin
              dma2mem[39][15].run()  ;
            end

            begin
              gen[39][16].run()  ;
            end
            begin
              drv[39][16].run()  ;
            end
            begin
              dma2mem[39][16].run()  ;
            end

            begin
              gen[39][17].run()  ;
            end
            begin
              drv[39][17].run()  ;
            end
            begin
              dma2mem[39][17].run()  ;
            end

            begin
              gen[39][18].run()  ;
            end
            begin
              drv[39][18].run()  ;
            end
            begin
              dma2mem[39][18].run()  ;
            end

            begin
              gen[39][19].run()  ;
            end
            begin
              drv[39][19].run()  ;
            end
            begin
              dma2mem[39][19].run()  ;
            end

            begin
              gen[39][20].run()  ;
            end
            begin
              drv[39][20].run()  ;
            end
            begin
              dma2mem[39][20].run()  ;
            end

            begin
              gen[39][21].run()  ;
            end
            begin
              drv[39][21].run()  ;
            end
            begin
              dma2mem[39][21].run()  ;
            end

            begin
              gen[39][22].run()  ;
            end
            begin
              drv[39][22].run()  ;
            end
            begin
              dma2mem[39][22].run()  ;
            end

            begin
              gen[39][23].run()  ;
            end
            begin
              drv[39][23].run()  ;
            end
            begin
              dma2mem[39][23].run()  ;
            end

            begin
              gen[39][24].run()  ;
            end
            begin
              drv[39][24].run()  ;
            end
            begin
              dma2mem[39][24].run()  ;
            end

            begin
              gen[39][25].run()  ;
            end
            begin
              drv[39][25].run()  ;
            end
            begin
              dma2mem[39][25].run()  ;
            end

            begin
              gen[39][26].run()  ;
            end
            begin
              drv[39][26].run()  ;
            end
            begin
              dma2mem[39][26].run()  ;
            end

            begin
              gen[39][27].run()  ;
            end
            begin
              drv[39][27].run()  ;
            end
            begin
              dma2mem[39][27].run()  ;
            end

            begin
              gen[39][28].run()  ;
            end
            begin
              drv[39][28].run()  ;
            end
            begin
              dma2mem[39][28].run()  ;
            end

            begin
              gen[39][29].run()  ;
            end
            begin
              drv[39][29].run()  ;
            end
            begin
              dma2mem[39][29].run()  ;
            end

            begin
              gen[39][30].run()  ;
            end
            begin
              drv[39][30].run()  ;
            end
            begin
              dma2mem[39][30].run()  ;
            end

            begin
              gen[39][31].run()  ;
            end
            begin
              drv[39][31].run()  ;
            end
            begin
              dma2mem[39][31].run()  ;
            end

            begin
              gen[40][0].run()  ;
            end
            begin
              drv[40][0].run()  ;
            end
            begin
              dma2mem[40][0].run()  ;
            end

            begin
              gen[40][1].run()  ;
            end
            begin
              drv[40][1].run()  ;
            end
            begin
              dma2mem[40][1].run()  ;
            end

            begin
              gen[40][2].run()  ;
            end
            begin
              drv[40][2].run()  ;
            end
            begin
              dma2mem[40][2].run()  ;
            end

            begin
              gen[40][3].run()  ;
            end
            begin
              drv[40][3].run()  ;
            end
            begin
              dma2mem[40][3].run()  ;
            end

            begin
              gen[40][4].run()  ;
            end
            begin
              drv[40][4].run()  ;
            end
            begin
              dma2mem[40][4].run()  ;
            end

            begin
              gen[40][5].run()  ;
            end
            begin
              drv[40][5].run()  ;
            end
            begin
              dma2mem[40][5].run()  ;
            end

            begin
              gen[40][6].run()  ;
            end
            begin
              drv[40][6].run()  ;
            end
            begin
              dma2mem[40][6].run()  ;
            end

            begin
              gen[40][7].run()  ;
            end
            begin
              drv[40][7].run()  ;
            end
            begin
              dma2mem[40][7].run()  ;
            end

            begin
              gen[40][8].run()  ;
            end
            begin
              drv[40][8].run()  ;
            end
            begin
              dma2mem[40][8].run()  ;
            end

            begin
              gen[40][9].run()  ;
            end
            begin
              drv[40][9].run()  ;
            end
            begin
              dma2mem[40][9].run()  ;
            end

            begin
              gen[40][10].run()  ;
            end
            begin
              drv[40][10].run()  ;
            end
            begin
              dma2mem[40][10].run()  ;
            end

            begin
              gen[40][11].run()  ;
            end
            begin
              drv[40][11].run()  ;
            end
            begin
              dma2mem[40][11].run()  ;
            end

            begin
              gen[40][12].run()  ;
            end
            begin
              drv[40][12].run()  ;
            end
            begin
              dma2mem[40][12].run()  ;
            end

            begin
              gen[40][13].run()  ;
            end
            begin
              drv[40][13].run()  ;
            end
            begin
              dma2mem[40][13].run()  ;
            end

            begin
              gen[40][14].run()  ;
            end
            begin
              drv[40][14].run()  ;
            end
            begin
              dma2mem[40][14].run()  ;
            end

            begin
              gen[40][15].run()  ;
            end
            begin
              drv[40][15].run()  ;
            end
            begin
              dma2mem[40][15].run()  ;
            end

            begin
              gen[40][16].run()  ;
            end
            begin
              drv[40][16].run()  ;
            end
            begin
              dma2mem[40][16].run()  ;
            end

            begin
              gen[40][17].run()  ;
            end
            begin
              drv[40][17].run()  ;
            end
            begin
              dma2mem[40][17].run()  ;
            end

            begin
              gen[40][18].run()  ;
            end
            begin
              drv[40][18].run()  ;
            end
            begin
              dma2mem[40][18].run()  ;
            end

            begin
              gen[40][19].run()  ;
            end
            begin
              drv[40][19].run()  ;
            end
            begin
              dma2mem[40][19].run()  ;
            end

            begin
              gen[40][20].run()  ;
            end
            begin
              drv[40][20].run()  ;
            end
            begin
              dma2mem[40][20].run()  ;
            end

            begin
              gen[40][21].run()  ;
            end
            begin
              drv[40][21].run()  ;
            end
            begin
              dma2mem[40][21].run()  ;
            end

            begin
              gen[40][22].run()  ;
            end
            begin
              drv[40][22].run()  ;
            end
            begin
              dma2mem[40][22].run()  ;
            end

            begin
              gen[40][23].run()  ;
            end
            begin
              drv[40][23].run()  ;
            end
            begin
              dma2mem[40][23].run()  ;
            end

            begin
              gen[40][24].run()  ;
            end
            begin
              drv[40][24].run()  ;
            end
            begin
              dma2mem[40][24].run()  ;
            end

            begin
              gen[40][25].run()  ;
            end
            begin
              drv[40][25].run()  ;
            end
            begin
              dma2mem[40][25].run()  ;
            end

            begin
              gen[40][26].run()  ;
            end
            begin
              drv[40][26].run()  ;
            end
            begin
              dma2mem[40][26].run()  ;
            end

            begin
              gen[40][27].run()  ;
            end
            begin
              drv[40][27].run()  ;
            end
            begin
              dma2mem[40][27].run()  ;
            end

            begin
              gen[40][28].run()  ;
            end
            begin
              drv[40][28].run()  ;
            end
            begin
              dma2mem[40][28].run()  ;
            end

            begin
              gen[40][29].run()  ;
            end
            begin
              drv[40][29].run()  ;
            end
            begin
              dma2mem[40][29].run()  ;
            end

            begin
              gen[40][30].run()  ;
            end
            begin
              drv[40][30].run()  ;
            end
            begin
              dma2mem[40][30].run()  ;
            end

            begin
              gen[40][31].run()  ;
            end
            begin
              drv[40][31].run()  ;
            end
            begin
              dma2mem[40][31].run()  ;
            end

            begin
              gen[41][0].run()  ;
            end
            begin
              drv[41][0].run()  ;
            end
            begin
              dma2mem[41][0].run()  ;
            end

            begin
              gen[41][1].run()  ;
            end
            begin
              drv[41][1].run()  ;
            end
            begin
              dma2mem[41][1].run()  ;
            end

            begin
              gen[41][2].run()  ;
            end
            begin
              drv[41][2].run()  ;
            end
            begin
              dma2mem[41][2].run()  ;
            end

            begin
              gen[41][3].run()  ;
            end
            begin
              drv[41][3].run()  ;
            end
            begin
              dma2mem[41][3].run()  ;
            end

            begin
              gen[41][4].run()  ;
            end
            begin
              drv[41][4].run()  ;
            end
            begin
              dma2mem[41][4].run()  ;
            end

            begin
              gen[41][5].run()  ;
            end
            begin
              drv[41][5].run()  ;
            end
            begin
              dma2mem[41][5].run()  ;
            end

            begin
              gen[41][6].run()  ;
            end
            begin
              drv[41][6].run()  ;
            end
            begin
              dma2mem[41][6].run()  ;
            end

            begin
              gen[41][7].run()  ;
            end
            begin
              drv[41][7].run()  ;
            end
            begin
              dma2mem[41][7].run()  ;
            end

            begin
              gen[41][8].run()  ;
            end
            begin
              drv[41][8].run()  ;
            end
            begin
              dma2mem[41][8].run()  ;
            end

            begin
              gen[41][9].run()  ;
            end
            begin
              drv[41][9].run()  ;
            end
            begin
              dma2mem[41][9].run()  ;
            end

            begin
              gen[41][10].run()  ;
            end
            begin
              drv[41][10].run()  ;
            end
            begin
              dma2mem[41][10].run()  ;
            end

            begin
              gen[41][11].run()  ;
            end
            begin
              drv[41][11].run()  ;
            end
            begin
              dma2mem[41][11].run()  ;
            end

            begin
              gen[41][12].run()  ;
            end
            begin
              drv[41][12].run()  ;
            end
            begin
              dma2mem[41][12].run()  ;
            end

            begin
              gen[41][13].run()  ;
            end
            begin
              drv[41][13].run()  ;
            end
            begin
              dma2mem[41][13].run()  ;
            end

            begin
              gen[41][14].run()  ;
            end
            begin
              drv[41][14].run()  ;
            end
            begin
              dma2mem[41][14].run()  ;
            end

            begin
              gen[41][15].run()  ;
            end
            begin
              drv[41][15].run()  ;
            end
            begin
              dma2mem[41][15].run()  ;
            end

            begin
              gen[41][16].run()  ;
            end
            begin
              drv[41][16].run()  ;
            end
            begin
              dma2mem[41][16].run()  ;
            end

            begin
              gen[41][17].run()  ;
            end
            begin
              drv[41][17].run()  ;
            end
            begin
              dma2mem[41][17].run()  ;
            end

            begin
              gen[41][18].run()  ;
            end
            begin
              drv[41][18].run()  ;
            end
            begin
              dma2mem[41][18].run()  ;
            end

            begin
              gen[41][19].run()  ;
            end
            begin
              drv[41][19].run()  ;
            end
            begin
              dma2mem[41][19].run()  ;
            end

            begin
              gen[41][20].run()  ;
            end
            begin
              drv[41][20].run()  ;
            end
            begin
              dma2mem[41][20].run()  ;
            end

            begin
              gen[41][21].run()  ;
            end
            begin
              drv[41][21].run()  ;
            end
            begin
              dma2mem[41][21].run()  ;
            end

            begin
              gen[41][22].run()  ;
            end
            begin
              drv[41][22].run()  ;
            end
            begin
              dma2mem[41][22].run()  ;
            end

            begin
              gen[41][23].run()  ;
            end
            begin
              drv[41][23].run()  ;
            end
            begin
              dma2mem[41][23].run()  ;
            end

            begin
              gen[41][24].run()  ;
            end
            begin
              drv[41][24].run()  ;
            end
            begin
              dma2mem[41][24].run()  ;
            end

            begin
              gen[41][25].run()  ;
            end
            begin
              drv[41][25].run()  ;
            end
            begin
              dma2mem[41][25].run()  ;
            end

            begin
              gen[41][26].run()  ;
            end
            begin
              drv[41][26].run()  ;
            end
            begin
              dma2mem[41][26].run()  ;
            end

            begin
              gen[41][27].run()  ;
            end
            begin
              drv[41][27].run()  ;
            end
            begin
              dma2mem[41][27].run()  ;
            end

            begin
              gen[41][28].run()  ;
            end
            begin
              drv[41][28].run()  ;
            end
            begin
              dma2mem[41][28].run()  ;
            end

            begin
              gen[41][29].run()  ;
            end
            begin
              drv[41][29].run()  ;
            end
            begin
              dma2mem[41][29].run()  ;
            end

            begin
              gen[41][30].run()  ;
            end
            begin
              drv[41][30].run()  ;
            end
            begin
              dma2mem[41][30].run()  ;
            end

            begin
              gen[41][31].run()  ;
            end
            begin
              drv[41][31].run()  ;
            end
            begin
              dma2mem[41][31].run()  ;
            end

            begin
              gen[42][0].run()  ;
            end
            begin
              drv[42][0].run()  ;
            end
            begin
              dma2mem[42][0].run()  ;
            end

            begin
              gen[42][1].run()  ;
            end
            begin
              drv[42][1].run()  ;
            end
            begin
              dma2mem[42][1].run()  ;
            end

            begin
              gen[42][2].run()  ;
            end
            begin
              drv[42][2].run()  ;
            end
            begin
              dma2mem[42][2].run()  ;
            end

            begin
              gen[42][3].run()  ;
            end
            begin
              drv[42][3].run()  ;
            end
            begin
              dma2mem[42][3].run()  ;
            end

            begin
              gen[42][4].run()  ;
            end
            begin
              drv[42][4].run()  ;
            end
            begin
              dma2mem[42][4].run()  ;
            end

            begin
              gen[42][5].run()  ;
            end
            begin
              drv[42][5].run()  ;
            end
            begin
              dma2mem[42][5].run()  ;
            end

            begin
              gen[42][6].run()  ;
            end
            begin
              drv[42][6].run()  ;
            end
            begin
              dma2mem[42][6].run()  ;
            end

            begin
              gen[42][7].run()  ;
            end
            begin
              drv[42][7].run()  ;
            end
            begin
              dma2mem[42][7].run()  ;
            end

            begin
              gen[42][8].run()  ;
            end
            begin
              drv[42][8].run()  ;
            end
            begin
              dma2mem[42][8].run()  ;
            end

            begin
              gen[42][9].run()  ;
            end
            begin
              drv[42][9].run()  ;
            end
            begin
              dma2mem[42][9].run()  ;
            end

            begin
              gen[42][10].run()  ;
            end
            begin
              drv[42][10].run()  ;
            end
            begin
              dma2mem[42][10].run()  ;
            end

            begin
              gen[42][11].run()  ;
            end
            begin
              drv[42][11].run()  ;
            end
            begin
              dma2mem[42][11].run()  ;
            end

            begin
              gen[42][12].run()  ;
            end
            begin
              drv[42][12].run()  ;
            end
            begin
              dma2mem[42][12].run()  ;
            end

            begin
              gen[42][13].run()  ;
            end
            begin
              drv[42][13].run()  ;
            end
            begin
              dma2mem[42][13].run()  ;
            end

            begin
              gen[42][14].run()  ;
            end
            begin
              drv[42][14].run()  ;
            end
            begin
              dma2mem[42][14].run()  ;
            end

            begin
              gen[42][15].run()  ;
            end
            begin
              drv[42][15].run()  ;
            end
            begin
              dma2mem[42][15].run()  ;
            end

            begin
              gen[42][16].run()  ;
            end
            begin
              drv[42][16].run()  ;
            end
            begin
              dma2mem[42][16].run()  ;
            end

            begin
              gen[42][17].run()  ;
            end
            begin
              drv[42][17].run()  ;
            end
            begin
              dma2mem[42][17].run()  ;
            end

            begin
              gen[42][18].run()  ;
            end
            begin
              drv[42][18].run()  ;
            end
            begin
              dma2mem[42][18].run()  ;
            end

            begin
              gen[42][19].run()  ;
            end
            begin
              drv[42][19].run()  ;
            end
            begin
              dma2mem[42][19].run()  ;
            end

            begin
              gen[42][20].run()  ;
            end
            begin
              drv[42][20].run()  ;
            end
            begin
              dma2mem[42][20].run()  ;
            end

            begin
              gen[42][21].run()  ;
            end
            begin
              drv[42][21].run()  ;
            end
            begin
              dma2mem[42][21].run()  ;
            end

            begin
              gen[42][22].run()  ;
            end
            begin
              drv[42][22].run()  ;
            end
            begin
              dma2mem[42][22].run()  ;
            end

            begin
              gen[42][23].run()  ;
            end
            begin
              drv[42][23].run()  ;
            end
            begin
              dma2mem[42][23].run()  ;
            end

            begin
              gen[42][24].run()  ;
            end
            begin
              drv[42][24].run()  ;
            end
            begin
              dma2mem[42][24].run()  ;
            end

            begin
              gen[42][25].run()  ;
            end
            begin
              drv[42][25].run()  ;
            end
            begin
              dma2mem[42][25].run()  ;
            end

            begin
              gen[42][26].run()  ;
            end
            begin
              drv[42][26].run()  ;
            end
            begin
              dma2mem[42][26].run()  ;
            end

            begin
              gen[42][27].run()  ;
            end
            begin
              drv[42][27].run()  ;
            end
            begin
              dma2mem[42][27].run()  ;
            end

            begin
              gen[42][28].run()  ;
            end
            begin
              drv[42][28].run()  ;
            end
            begin
              dma2mem[42][28].run()  ;
            end

            begin
              gen[42][29].run()  ;
            end
            begin
              drv[42][29].run()  ;
            end
            begin
              dma2mem[42][29].run()  ;
            end

            begin
              gen[42][30].run()  ;
            end
            begin
              drv[42][30].run()  ;
            end
            begin
              dma2mem[42][30].run()  ;
            end

            begin
              gen[42][31].run()  ;
            end
            begin
              drv[42][31].run()  ;
            end
            begin
              dma2mem[42][31].run()  ;
            end

            begin
              gen[43][0].run()  ;
            end
            begin
              drv[43][0].run()  ;
            end
            begin
              dma2mem[43][0].run()  ;
            end

            begin
              gen[43][1].run()  ;
            end
            begin
              drv[43][1].run()  ;
            end
            begin
              dma2mem[43][1].run()  ;
            end

            begin
              gen[43][2].run()  ;
            end
            begin
              drv[43][2].run()  ;
            end
            begin
              dma2mem[43][2].run()  ;
            end

            begin
              gen[43][3].run()  ;
            end
            begin
              drv[43][3].run()  ;
            end
            begin
              dma2mem[43][3].run()  ;
            end

            begin
              gen[43][4].run()  ;
            end
            begin
              drv[43][4].run()  ;
            end
            begin
              dma2mem[43][4].run()  ;
            end

            begin
              gen[43][5].run()  ;
            end
            begin
              drv[43][5].run()  ;
            end
            begin
              dma2mem[43][5].run()  ;
            end

            begin
              gen[43][6].run()  ;
            end
            begin
              drv[43][6].run()  ;
            end
            begin
              dma2mem[43][6].run()  ;
            end

            begin
              gen[43][7].run()  ;
            end
            begin
              drv[43][7].run()  ;
            end
            begin
              dma2mem[43][7].run()  ;
            end

            begin
              gen[43][8].run()  ;
            end
            begin
              drv[43][8].run()  ;
            end
            begin
              dma2mem[43][8].run()  ;
            end

            begin
              gen[43][9].run()  ;
            end
            begin
              drv[43][9].run()  ;
            end
            begin
              dma2mem[43][9].run()  ;
            end

            begin
              gen[43][10].run()  ;
            end
            begin
              drv[43][10].run()  ;
            end
            begin
              dma2mem[43][10].run()  ;
            end

            begin
              gen[43][11].run()  ;
            end
            begin
              drv[43][11].run()  ;
            end
            begin
              dma2mem[43][11].run()  ;
            end

            begin
              gen[43][12].run()  ;
            end
            begin
              drv[43][12].run()  ;
            end
            begin
              dma2mem[43][12].run()  ;
            end

            begin
              gen[43][13].run()  ;
            end
            begin
              drv[43][13].run()  ;
            end
            begin
              dma2mem[43][13].run()  ;
            end

            begin
              gen[43][14].run()  ;
            end
            begin
              drv[43][14].run()  ;
            end
            begin
              dma2mem[43][14].run()  ;
            end

            begin
              gen[43][15].run()  ;
            end
            begin
              drv[43][15].run()  ;
            end
            begin
              dma2mem[43][15].run()  ;
            end

            begin
              gen[43][16].run()  ;
            end
            begin
              drv[43][16].run()  ;
            end
            begin
              dma2mem[43][16].run()  ;
            end

            begin
              gen[43][17].run()  ;
            end
            begin
              drv[43][17].run()  ;
            end
            begin
              dma2mem[43][17].run()  ;
            end

            begin
              gen[43][18].run()  ;
            end
            begin
              drv[43][18].run()  ;
            end
            begin
              dma2mem[43][18].run()  ;
            end

            begin
              gen[43][19].run()  ;
            end
            begin
              drv[43][19].run()  ;
            end
            begin
              dma2mem[43][19].run()  ;
            end

            begin
              gen[43][20].run()  ;
            end
            begin
              drv[43][20].run()  ;
            end
            begin
              dma2mem[43][20].run()  ;
            end

            begin
              gen[43][21].run()  ;
            end
            begin
              drv[43][21].run()  ;
            end
            begin
              dma2mem[43][21].run()  ;
            end

            begin
              gen[43][22].run()  ;
            end
            begin
              drv[43][22].run()  ;
            end
            begin
              dma2mem[43][22].run()  ;
            end

            begin
              gen[43][23].run()  ;
            end
            begin
              drv[43][23].run()  ;
            end
            begin
              dma2mem[43][23].run()  ;
            end

            begin
              gen[43][24].run()  ;
            end
            begin
              drv[43][24].run()  ;
            end
            begin
              dma2mem[43][24].run()  ;
            end

            begin
              gen[43][25].run()  ;
            end
            begin
              drv[43][25].run()  ;
            end
            begin
              dma2mem[43][25].run()  ;
            end

            begin
              gen[43][26].run()  ;
            end
            begin
              drv[43][26].run()  ;
            end
            begin
              dma2mem[43][26].run()  ;
            end

            begin
              gen[43][27].run()  ;
            end
            begin
              drv[43][27].run()  ;
            end
            begin
              dma2mem[43][27].run()  ;
            end

            begin
              gen[43][28].run()  ;
            end
            begin
              drv[43][28].run()  ;
            end
            begin
              dma2mem[43][28].run()  ;
            end

            begin
              gen[43][29].run()  ;
            end
            begin
              drv[43][29].run()  ;
            end
            begin
              dma2mem[43][29].run()  ;
            end

            begin
              gen[43][30].run()  ;
            end
            begin
              drv[43][30].run()  ;
            end
            begin
              dma2mem[43][30].run()  ;
            end

            begin
              gen[43][31].run()  ;
            end
            begin
              drv[43][31].run()  ;
            end
            begin
              dma2mem[43][31].run()  ;
            end

            begin
              gen[44][0].run()  ;
            end
            begin
              drv[44][0].run()  ;
            end
            begin
              dma2mem[44][0].run()  ;
            end

            begin
              gen[44][1].run()  ;
            end
            begin
              drv[44][1].run()  ;
            end
            begin
              dma2mem[44][1].run()  ;
            end

            begin
              gen[44][2].run()  ;
            end
            begin
              drv[44][2].run()  ;
            end
            begin
              dma2mem[44][2].run()  ;
            end

            begin
              gen[44][3].run()  ;
            end
            begin
              drv[44][3].run()  ;
            end
            begin
              dma2mem[44][3].run()  ;
            end

            begin
              gen[44][4].run()  ;
            end
            begin
              drv[44][4].run()  ;
            end
            begin
              dma2mem[44][4].run()  ;
            end

            begin
              gen[44][5].run()  ;
            end
            begin
              drv[44][5].run()  ;
            end
            begin
              dma2mem[44][5].run()  ;
            end

            begin
              gen[44][6].run()  ;
            end
            begin
              drv[44][6].run()  ;
            end
            begin
              dma2mem[44][6].run()  ;
            end

            begin
              gen[44][7].run()  ;
            end
            begin
              drv[44][7].run()  ;
            end
            begin
              dma2mem[44][7].run()  ;
            end

            begin
              gen[44][8].run()  ;
            end
            begin
              drv[44][8].run()  ;
            end
            begin
              dma2mem[44][8].run()  ;
            end

            begin
              gen[44][9].run()  ;
            end
            begin
              drv[44][9].run()  ;
            end
            begin
              dma2mem[44][9].run()  ;
            end

            begin
              gen[44][10].run()  ;
            end
            begin
              drv[44][10].run()  ;
            end
            begin
              dma2mem[44][10].run()  ;
            end

            begin
              gen[44][11].run()  ;
            end
            begin
              drv[44][11].run()  ;
            end
            begin
              dma2mem[44][11].run()  ;
            end

            begin
              gen[44][12].run()  ;
            end
            begin
              drv[44][12].run()  ;
            end
            begin
              dma2mem[44][12].run()  ;
            end

            begin
              gen[44][13].run()  ;
            end
            begin
              drv[44][13].run()  ;
            end
            begin
              dma2mem[44][13].run()  ;
            end

            begin
              gen[44][14].run()  ;
            end
            begin
              drv[44][14].run()  ;
            end
            begin
              dma2mem[44][14].run()  ;
            end

            begin
              gen[44][15].run()  ;
            end
            begin
              drv[44][15].run()  ;
            end
            begin
              dma2mem[44][15].run()  ;
            end

            begin
              gen[44][16].run()  ;
            end
            begin
              drv[44][16].run()  ;
            end
            begin
              dma2mem[44][16].run()  ;
            end

            begin
              gen[44][17].run()  ;
            end
            begin
              drv[44][17].run()  ;
            end
            begin
              dma2mem[44][17].run()  ;
            end

            begin
              gen[44][18].run()  ;
            end
            begin
              drv[44][18].run()  ;
            end
            begin
              dma2mem[44][18].run()  ;
            end

            begin
              gen[44][19].run()  ;
            end
            begin
              drv[44][19].run()  ;
            end
            begin
              dma2mem[44][19].run()  ;
            end

            begin
              gen[44][20].run()  ;
            end
            begin
              drv[44][20].run()  ;
            end
            begin
              dma2mem[44][20].run()  ;
            end

            begin
              gen[44][21].run()  ;
            end
            begin
              drv[44][21].run()  ;
            end
            begin
              dma2mem[44][21].run()  ;
            end

            begin
              gen[44][22].run()  ;
            end
            begin
              drv[44][22].run()  ;
            end
            begin
              dma2mem[44][22].run()  ;
            end

            begin
              gen[44][23].run()  ;
            end
            begin
              drv[44][23].run()  ;
            end
            begin
              dma2mem[44][23].run()  ;
            end

            begin
              gen[44][24].run()  ;
            end
            begin
              drv[44][24].run()  ;
            end
            begin
              dma2mem[44][24].run()  ;
            end

            begin
              gen[44][25].run()  ;
            end
            begin
              drv[44][25].run()  ;
            end
            begin
              dma2mem[44][25].run()  ;
            end

            begin
              gen[44][26].run()  ;
            end
            begin
              drv[44][26].run()  ;
            end
            begin
              dma2mem[44][26].run()  ;
            end

            begin
              gen[44][27].run()  ;
            end
            begin
              drv[44][27].run()  ;
            end
            begin
              dma2mem[44][27].run()  ;
            end

            begin
              gen[44][28].run()  ;
            end
            begin
              drv[44][28].run()  ;
            end
            begin
              dma2mem[44][28].run()  ;
            end

            begin
              gen[44][29].run()  ;
            end
            begin
              drv[44][29].run()  ;
            end
            begin
              dma2mem[44][29].run()  ;
            end

            begin
              gen[44][30].run()  ;
            end
            begin
              drv[44][30].run()  ;
            end
            begin
              dma2mem[44][30].run()  ;
            end

            begin
              gen[44][31].run()  ;
            end
            begin
              drv[44][31].run()  ;
            end
            begin
              dma2mem[44][31].run()  ;
            end

            begin
              gen[45][0].run()  ;
            end
            begin
              drv[45][0].run()  ;
            end
            begin
              dma2mem[45][0].run()  ;
            end

            begin
              gen[45][1].run()  ;
            end
            begin
              drv[45][1].run()  ;
            end
            begin
              dma2mem[45][1].run()  ;
            end

            begin
              gen[45][2].run()  ;
            end
            begin
              drv[45][2].run()  ;
            end
            begin
              dma2mem[45][2].run()  ;
            end

            begin
              gen[45][3].run()  ;
            end
            begin
              drv[45][3].run()  ;
            end
            begin
              dma2mem[45][3].run()  ;
            end

            begin
              gen[45][4].run()  ;
            end
            begin
              drv[45][4].run()  ;
            end
            begin
              dma2mem[45][4].run()  ;
            end

            begin
              gen[45][5].run()  ;
            end
            begin
              drv[45][5].run()  ;
            end
            begin
              dma2mem[45][5].run()  ;
            end

            begin
              gen[45][6].run()  ;
            end
            begin
              drv[45][6].run()  ;
            end
            begin
              dma2mem[45][6].run()  ;
            end

            begin
              gen[45][7].run()  ;
            end
            begin
              drv[45][7].run()  ;
            end
            begin
              dma2mem[45][7].run()  ;
            end

            begin
              gen[45][8].run()  ;
            end
            begin
              drv[45][8].run()  ;
            end
            begin
              dma2mem[45][8].run()  ;
            end

            begin
              gen[45][9].run()  ;
            end
            begin
              drv[45][9].run()  ;
            end
            begin
              dma2mem[45][9].run()  ;
            end

            begin
              gen[45][10].run()  ;
            end
            begin
              drv[45][10].run()  ;
            end
            begin
              dma2mem[45][10].run()  ;
            end

            begin
              gen[45][11].run()  ;
            end
            begin
              drv[45][11].run()  ;
            end
            begin
              dma2mem[45][11].run()  ;
            end

            begin
              gen[45][12].run()  ;
            end
            begin
              drv[45][12].run()  ;
            end
            begin
              dma2mem[45][12].run()  ;
            end

            begin
              gen[45][13].run()  ;
            end
            begin
              drv[45][13].run()  ;
            end
            begin
              dma2mem[45][13].run()  ;
            end

            begin
              gen[45][14].run()  ;
            end
            begin
              drv[45][14].run()  ;
            end
            begin
              dma2mem[45][14].run()  ;
            end

            begin
              gen[45][15].run()  ;
            end
            begin
              drv[45][15].run()  ;
            end
            begin
              dma2mem[45][15].run()  ;
            end

            begin
              gen[45][16].run()  ;
            end
            begin
              drv[45][16].run()  ;
            end
            begin
              dma2mem[45][16].run()  ;
            end

            begin
              gen[45][17].run()  ;
            end
            begin
              drv[45][17].run()  ;
            end
            begin
              dma2mem[45][17].run()  ;
            end

            begin
              gen[45][18].run()  ;
            end
            begin
              drv[45][18].run()  ;
            end
            begin
              dma2mem[45][18].run()  ;
            end

            begin
              gen[45][19].run()  ;
            end
            begin
              drv[45][19].run()  ;
            end
            begin
              dma2mem[45][19].run()  ;
            end

            begin
              gen[45][20].run()  ;
            end
            begin
              drv[45][20].run()  ;
            end
            begin
              dma2mem[45][20].run()  ;
            end

            begin
              gen[45][21].run()  ;
            end
            begin
              drv[45][21].run()  ;
            end
            begin
              dma2mem[45][21].run()  ;
            end

            begin
              gen[45][22].run()  ;
            end
            begin
              drv[45][22].run()  ;
            end
            begin
              dma2mem[45][22].run()  ;
            end

            begin
              gen[45][23].run()  ;
            end
            begin
              drv[45][23].run()  ;
            end
            begin
              dma2mem[45][23].run()  ;
            end

            begin
              gen[45][24].run()  ;
            end
            begin
              drv[45][24].run()  ;
            end
            begin
              dma2mem[45][24].run()  ;
            end

            begin
              gen[45][25].run()  ;
            end
            begin
              drv[45][25].run()  ;
            end
            begin
              dma2mem[45][25].run()  ;
            end

            begin
              gen[45][26].run()  ;
            end
            begin
              drv[45][26].run()  ;
            end
            begin
              dma2mem[45][26].run()  ;
            end

            begin
              gen[45][27].run()  ;
            end
            begin
              drv[45][27].run()  ;
            end
            begin
              dma2mem[45][27].run()  ;
            end

            begin
              gen[45][28].run()  ;
            end
            begin
              drv[45][28].run()  ;
            end
            begin
              dma2mem[45][28].run()  ;
            end

            begin
              gen[45][29].run()  ;
            end
            begin
              drv[45][29].run()  ;
            end
            begin
              dma2mem[45][29].run()  ;
            end

            begin
              gen[45][30].run()  ;
            end
            begin
              drv[45][30].run()  ;
            end
            begin
              dma2mem[45][30].run()  ;
            end

            begin
              gen[45][31].run()  ;
            end
            begin
              drv[45][31].run()  ;
            end
            begin
              dma2mem[45][31].run()  ;
            end

            begin
              gen[46][0].run()  ;
            end
            begin
              drv[46][0].run()  ;
            end
            begin
              dma2mem[46][0].run()  ;
            end

            begin
              gen[46][1].run()  ;
            end
            begin
              drv[46][1].run()  ;
            end
            begin
              dma2mem[46][1].run()  ;
            end

            begin
              gen[46][2].run()  ;
            end
            begin
              drv[46][2].run()  ;
            end
            begin
              dma2mem[46][2].run()  ;
            end

            begin
              gen[46][3].run()  ;
            end
            begin
              drv[46][3].run()  ;
            end
            begin
              dma2mem[46][3].run()  ;
            end

            begin
              gen[46][4].run()  ;
            end
            begin
              drv[46][4].run()  ;
            end
            begin
              dma2mem[46][4].run()  ;
            end

            begin
              gen[46][5].run()  ;
            end
            begin
              drv[46][5].run()  ;
            end
            begin
              dma2mem[46][5].run()  ;
            end

            begin
              gen[46][6].run()  ;
            end
            begin
              drv[46][6].run()  ;
            end
            begin
              dma2mem[46][6].run()  ;
            end

            begin
              gen[46][7].run()  ;
            end
            begin
              drv[46][7].run()  ;
            end
            begin
              dma2mem[46][7].run()  ;
            end

            begin
              gen[46][8].run()  ;
            end
            begin
              drv[46][8].run()  ;
            end
            begin
              dma2mem[46][8].run()  ;
            end

            begin
              gen[46][9].run()  ;
            end
            begin
              drv[46][9].run()  ;
            end
            begin
              dma2mem[46][9].run()  ;
            end

            begin
              gen[46][10].run()  ;
            end
            begin
              drv[46][10].run()  ;
            end
            begin
              dma2mem[46][10].run()  ;
            end

            begin
              gen[46][11].run()  ;
            end
            begin
              drv[46][11].run()  ;
            end
            begin
              dma2mem[46][11].run()  ;
            end

            begin
              gen[46][12].run()  ;
            end
            begin
              drv[46][12].run()  ;
            end
            begin
              dma2mem[46][12].run()  ;
            end

            begin
              gen[46][13].run()  ;
            end
            begin
              drv[46][13].run()  ;
            end
            begin
              dma2mem[46][13].run()  ;
            end

            begin
              gen[46][14].run()  ;
            end
            begin
              drv[46][14].run()  ;
            end
            begin
              dma2mem[46][14].run()  ;
            end

            begin
              gen[46][15].run()  ;
            end
            begin
              drv[46][15].run()  ;
            end
            begin
              dma2mem[46][15].run()  ;
            end

            begin
              gen[46][16].run()  ;
            end
            begin
              drv[46][16].run()  ;
            end
            begin
              dma2mem[46][16].run()  ;
            end

            begin
              gen[46][17].run()  ;
            end
            begin
              drv[46][17].run()  ;
            end
            begin
              dma2mem[46][17].run()  ;
            end

            begin
              gen[46][18].run()  ;
            end
            begin
              drv[46][18].run()  ;
            end
            begin
              dma2mem[46][18].run()  ;
            end

            begin
              gen[46][19].run()  ;
            end
            begin
              drv[46][19].run()  ;
            end
            begin
              dma2mem[46][19].run()  ;
            end

            begin
              gen[46][20].run()  ;
            end
            begin
              drv[46][20].run()  ;
            end
            begin
              dma2mem[46][20].run()  ;
            end

            begin
              gen[46][21].run()  ;
            end
            begin
              drv[46][21].run()  ;
            end
            begin
              dma2mem[46][21].run()  ;
            end

            begin
              gen[46][22].run()  ;
            end
            begin
              drv[46][22].run()  ;
            end
            begin
              dma2mem[46][22].run()  ;
            end

            begin
              gen[46][23].run()  ;
            end
            begin
              drv[46][23].run()  ;
            end
            begin
              dma2mem[46][23].run()  ;
            end

            begin
              gen[46][24].run()  ;
            end
            begin
              drv[46][24].run()  ;
            end
            begin
              dma2mem[46][24].run()  ;
            end

            begin
              gen[46][25].run()  ;
            end
            begin
              drv[46][25].run()  ;
            end
            begin
              dma2mem[46][25].run()  ;
            end

            begin
              gen[46][26].run()  ;
            end
            begin
              drv[46][26].run()  ;
            end
            begin
              dma2mem[46][26].run()  ;
            end

            begin
              gen[46][27].run()  ;
            end
            begin
              drv[46][27].run()  ;
            end
            begin
              dma2mem[46][27].run()  ;
            end

            begin
              gen[46][28].run()  ;
            end
            begin
              drv[46][28].run()  ;
            end
            begin
              dma2mem[46][28].run()  ;
            end

            begin
              gen[46][29].run()  ;
            end
            begin
              drv[46][29].run()  ;
            end
            begin
              dma2mem[46][29].run()  ;
            end

            begin
              gen[46][30].run()  ;
            end
            begin
              drv[46][30].run()  ;
            end
            begin
              dma2mem[46][30].run()  ;
            end

            begin
              gen[46][31].run()  ;
            end
            begin
              drv[46][31].run()  ;
            end
            begin
              dma2mem[46][31].run()  ;
            end

            begin
              gen[47][0].run()  ;
            end
            begin
              drv[47][0].run()  ;
            end
            begin
              dma2mem[47][0].run()  ;
            end

            begin
              gen[47][1].run()  ;
            end
            begin
              drv[47][1].run()  ;
            end
            begin
              dma2mem[47][1].run()  ;
            end

            begin
              gen[47][2].run()  ;
            end
            begin
              drv[47][2].run()  ;
            end
            begin
              dma2mem[47][2].run()  ;
            end

            begin
              gen[47][3].run()  ;
            end
            begin
              drv[47][3].run()  ;
            end
            begin
              dma2mem[47][3].run()  ;
            end

            begin
              gen[47][4].run()  ;
            end
            begin
              drv[47][4].run()  ;
            end
            begin
              dma2mem[47][4].run()  ;
            end

            begin
              gen[47][5].run()  ;
            end
            begin
              drv[47][5].run()  ;
            end
            begin
              dma2mem[47][5].run()  ;
            end

            begin
              gen[47][6].run()  ;
            end
            begin
              drv[47][6].run()  ;
            end
            begin
              dma2mem[47][6].run()  ;
            end

            begin
              gen[47][7].run()  ;
            end
            begin
              drv[47][7].run()  ;
            end
            begin
              dma2mem[47][7].run()  ;
            end

            begin
              gen[47][8].run()  ;
            end
            begin
              drv[47][8].run()  ;
            end
            begin
              dma2mem[47][8].run()  ;
            end

            begin
              gen[47][9].run()  ;
            end
            begin
              drv[47][9].run()  ;
            end
            begin
              dma2mem[47][9].run()  ;
            end

            begin
              gen[47][10].run()  ;
            end
            begin
              drv[47][10].run()  ;
            end
            begin
              dma2mem[47][10].run()  ;
            end

            begin
              gen[47][11].run()  ;
            end
            begin
              drv[47][11].run()  ;
            end
            begin
              dma2mem[47][11].run()  ;
            end

            begin
              gen[47][12].run()  ;
            end
            begin
              drv[47][12].run()  ;
            end
            begin
              dma2mem[47][12].run()  ;
            end

            begin
              gen[47][13].run()  ;
            end
            begin
              drv[47][13].run()  ;
            end
            begin
              dma2mem[47][13].run()  ;
            end

            begin
              gen[47][14].run()  ;
            end
            begin
              drv[47][14].run()  ;
            end
            begin
              dma2mem[47][14].run()  ;
            end

            begin
              gen[47][15].run()  ;
            end
            begin
              drv[47][15].run()  ;
            end
            begin
              dma2mem[47][15].run()  ;
            end

            begin
              gen[47][16].run()  ;
            end
            begin
              drv[47][16].run()  ;
            end
            begin
              dma2mem[47][16].run()  ;
            end

            begin
              gen[47][17].run()  ;
            end
            begin
              drv[47][17].run()  ;
            end
            begin
              dma2mem[47][17].run()  ;
            end

            begin
              gen[47][18].run()  ;
            end
            begin
              drv[47][18].run()  ;
            end
            begin
              dma2mem[47][18].run()  ;
            end

            begin
              gen[47][19].run()  ;
            end
            begin
              drv[47][19].run()  ;
            end
            begin
              dma2mem[47][19].run()  ;
            end

            begin
              gen[47][20].run()  ;
            end
            begin
              drv[47][20].run()  ;
            end
            begin
              dma2mem[47][20].run()  ;
            end

            begin
              gen[47][21].run()  ;
            end
            begin
              drv[47][21].run()  ;
            end
            begin
              dma2mem[47][21].run()  ;
            end

            begin
              gen[47][22].run()  ;
            end
            begin
              drv[47][22].run()  ;
            end
            begin
              dma2mem[47][22].run()  ;
            end

            begin
              gen[47][23].run()  ;
            end
            begin
              drv[47][23].run()  ;
            end
            begin
              dma2mem[47][23].run()  ;
            end

            begin
              gen[47][24].run()  ;
            end
            begin
              drv[47][24].run()  ;
            end
            begin
              dma2mem[47][24].run()  ;
            end

            begin
              gen[47][25].run()  ;
            end
            begin
              drv[47][25].run()  ;
            end
            begin
              dma2mem[47][25].run()  ;
            end

            begin
              gen[47][26].run()  ;
            end
            begin
              drv[47][26].run()  ;
            end
            begin
              dma2mem[47][26].run()  ;
            end

            begin
              gen[47][27].run()  ;
            end
            begin
              drv[47][27].run()  ;
            end
            begin
              dma2mem[47][27].run()  ;
            end

            begin
              gen[47][28].run()  ;
            end
            begin
              drv[47][28].run()  ;
            end
            begin
              dma2mem[47][28].run()  ;
            end

            begin
              gen[47][29].run()  ;
            end
            begin
              drv[47][29].run()  ;
            end
            begin
              dma2mem[47][29].run()  ;
            end

            begin
              gen[47][30].run()  ;
            end
            begin
              drv[47][30].run()  ;
            end
            begin
              dma2mem[47][30].run()  ;
            end

            begin
              gen[47][31].run()  ;
            end
            begin
              drv[47][31].run()  ;
            end
            begin
              dma2mem[47][31].run()  ;
            end

            begin
              gen[48][0].run()  ;
            end
            begin
              drv[48][0].run()  ;
            end
            begin
              dma2mem[48][0].run()  ;
            end

            begin
              gen[48][1].run()  ;
            end
            begin
              drv[48][1].run()  ;
            end
            begin
              dma2mem[48][1].run()  ;
            end

            begin
              gen[48][2].run()  ;
            end
            begin
              drv[48][2].run()  ;
            end
            begin
              dma2mem[48][2].run()  ;
            end

            begin
              gen[48][3].run()  ;
            end
            begin
              drv[48][3].run()  ;
            end
            begin
              dma2mem[48][3].run()  ;
            end

            begin
              gen[48][4].run()  ;
            end
            begin
              drv[48][4].run()  ;
            end
            begin
              dma2mem[48][4].run()  ;
            end

            begin
              gen[48][5].run()  ;
            end
            begin
              drv[48][5].run()  ;
            end
            begin
              dma2mem[48][5].run()  ;
            end

            begin
              gen[48][6].run()  ;
            end
            begin
              drv[48][6].run()  ;
            end
            begin
              dma2mem[48][6].run()  ;
            end

            begin
              gen[48][7].run()  ;
            end
            begin
              drv[48][7].run()  ;
            end
            begin
              dma2mem[48][7].run()  ;
            end

            begin
              gen[48][8].run()  ;
            end
            begin
              drv[48][8].run()  ;
            end
            begin
              dma2mem[48][8].run()  ;
            end

            begin
              gen[48][9].run()  ;
            end
            begin
              drv[48][9].run()  ;
            end
            begin
              dma2mem[48][9].run()  ;
            end

            begin
              gen[48][10].run()  ;
            end
            begin
              drv[48][10].run()  ;
            end
            begin
              dma2mem[48][10].run()  ;
            end

            begin
              gen[48][11].run()  ;
            end
            begin
              drv[48][11].run()  ;
            end
            begin
              dma2mem[48][11].run()  ;
            end

            begin
              gen[48][12].run()  ;
            end
            begin
              drv[48][12].run()  ;
            end
            begin
              dma2mem[48][12].run()  ;
            end

            begin
              gen[48][13].run()  ;
            end
            begin
              drv[48][13].run()  ;
            end
            begin
              dma2mem[48][13].run()  ;
            end

            begin
              gen[48][14].run()  ;
            end
            begin
              drv[48][14].run()  ;
            end
            begin
              dma2mem[48][14].run()  ;
            end

            begin
              gen[48][15].run()  ;
            end
            begin
              drv[48][15].run()  ;
            end
            begin
              dma2mem[48][15].run()  ;
            end

            begin
              gen[48][16].run()  ;
            end
            begin
              drv[48][16].run()  ;
            end
            begin
              dma2mem[48][16].run()  ;
            end

            begin
              gen[48][17].run()  ;
            end
            begin
              drv[48][17].run()  ;
            end
            begin
              dma2mem[48][17].run()  ;
            end

            begin
              gen[48][18].run()  ;
            end
            begin
              drv[48][18].run()  ;
            end
            begin
              dma2mem[48][18].run()  ;
            end

            begin
              gen[48][19].run()  ;
            end
            begin
              drv[48][19].run()  ;
            end
            begin
              dma2mem[48][19].run()  ;
            end

            begin
              gen[48][20].run()  ;
            end
            begin
              drv[48][20].run()  ;
            end
            begin
              dma2mem[48][20].run()  ;
            end

            begin
              gen[48][21].run()  ;
            end
            begin
              drv[48][21].run()  ;
            end
            begin
              dma2mem[48][21].run()  ;
            end

            begin
              gen[48][22].run()  ;
            end
            begin
              drv[48][22].run()  ;
            end
            begin
              dma2mem[48][22].run()  ;
            end

            begin
              gen[48][23].run()  ;
            end
            begin
              drv[48][23].run()  ;
            end
            begin
              dma2mem[48][23].run()  ;
            end

            begin
              gen[48][24].run()  ;
            end
            begin
              drv[48][24].run()  ;
            end
            begin
              dma2mem[48][24].run()  ;
            end

            begin
              gen[48][25].run()  ;
            end
            begin
              drv[48][25].run()  ;
            end
            begin
              dma2mem[48][25].run()  ;
            end

            begin
              gen[48][26].run()  ;
            end
            begin
              drv[48][26].run()  ;
            end
            begin
              dma2mem[48][26].run()  ;
            end

            begin
              gen[48][27].run()  ;
            end
            begin
              drv[48][27].run()  ;
            end
            begin
              dma2mem[48][27].run()  ;
            end

            begin
              gen[48][28].run()  ;
            end
            begin
              drv[48][28].run()  ;
            end
            begin
              dma2mem[48][28].run()  ;
            end

            begin
              gen[48][29].run()  ;
            end
            begin
              drv[48][29].run()  ;
            end
            begin
              dma2mem[48][29].run()  ;
            end

            begin
              gen[48][30].run()  ;
            end
            begin
              drv[48][30].run()  ;
            end
            begin
              dma2mem[48][30].run()  ;
            end

            begin
              gen[48][31].run()  ;
            end
            begin
              drv[48][31].run()  ;
            end
            begin
              dma2mem[48][31].run()  ;
            end

            begin
              gen[49][0].run()  ;
            end
            begin
              drv[49][0].run()  ;
            end
            begin
              dma2mem[49][0].run()  ;
            end

            begin
              gen[49][1].run()  ;
            end
            begin
              drv[49][1].run()  ;
            end
            begin
              dma2mem[49][1].run()  ;
            end

            begin
              gen[49][2].run()  ;
            end
            begin
              drv[49][2].run()  ;
            end
            begin
              dma2mem[49][2].run()  ;
            end

            begin
              gen[49][3].run()  ;
            end
            begin
              drv[49][3].run()  ;
            end
            begin
              dma2mem[49][3].run()  ;
            end

            begin
              gen[49][4].run()  ;
            end
            begin
              drv[49][4].run()  ;
            end
            begin
              dma2mem[49][4].run()  ;
            end

            begin
              gen[49][5].run()  ;
            end
            begin
              drv[49][5].run()  ;
            end
            begin
              dma2mem[49][5].run()  ;
            end

            begin
              gen[49][6].run()  ;
            end
            begin
              drv[49][6].run()  ;
            end
            begin
              dma2mem[49][6].run()  ;
            end

            begin
              gen[49][7].run()  ;
            end
            begin
              drv[49][7].run()  ;
            end
            begin
              dma2mem[49][7].run()  ;
            end

            begin
              gen[49][8].run()  ;
            end
            begin
              drv[49][8].run()  ;
            end
            begin
              dma2mem[49][8].run()  ;
            end

            begin
              gen[49][9].run()  ;
            end
            begin
              drv[49][9].run()  ;
            end
            begin
              dma2mem[49][9].run()  ;
            end

            begin
              gen[49][10].run()  ;
            end
            begin
              drv[49][10].run()  ;
            end
            begin
              dma2mem[49][10].run()  ;
            end

            begin
              gen[49][11].run()  ;
            end
            begin
              drv[49][11].run()  ;
            end
            begin
              dma2mem[49][11].run()  ;
            end

            begin
              gen[49][12].run()  ;
            end
            begin
              drv[49][12].run()  ;
            end
            begin
              dma2mem[49][12].run()  ;
            end

            begin
              gen[49][13].run()  ;
            end
            begin
              drv[49][13].run()  ;
            end
            begin
              dma2mem[49][13].run()  ;
            end

            begin
              gen[49][14].run()  ;
            end
            begin
              drv[49][14].run()  ;
            end
            begin
              dma2mem[49][14].run()  ;
            end

            begin
              gen[49][15].run()  ;
            end
            begin
              drv[49][15].run()  ;
            end
            begin
              dma2mem[49][15].run()  ;
            end

            begin
              gen[49][16].run()  ;
            end
            begin
              drv[49][16].run()  ;
            end
            begin
              dma2mem[49][16].run()  ;
            end

            begin
              gen[49][17].run()  ;
            end
            begin
              drv[49][17].run()  ;
            end
            begin
              dma2mem[49][17].run()  ;
            end

            begin
              gen[49][18].run()  ;
            end
            begin
              drv[49][18].run()  ;
            end
            begin
              dma2mem[49][18].run()  ;
            end

            begin
              gen[49][19].run()  ;
            end
            begin
              drv[49][19].run()  ;
            end
            begin
              dma2mem[49][19].run()  ;
            end

            begin
              gen[49][20].run()  ;
            end
            begin
              drv[49][20].run()  ;
            end
            begin
              dma2mem[49][20].run()  ;
            end

            begin
              gen[49][21].run()  ;
            end
            begin
              drv[49][21].run()  ;
            end
            begin
              dma2mem[49][21].run()  ;
            end

            begin
              gen[49][22].run()  ;
            end
            begin
              drv[49][22].run()  ;
            end
            begin
              dma2mem[49][22].run()  ;
            end

            begin
              gen[49][23].run()  ;
            end
            begin
              drv[49][23].run()  ;
            end
            begin
              dma2mem[49][23].run()  ;
            end

            begin
              gen[49][24].run()  ;
            end
            begin
              drv[49][24].run()  ;
            end
            begin
              dma2mem[49][24].run()  ;
            end

            begin
              gen[49][25].run()  ;
            end
            begin
              drv[49][25].run()  ;
            end
            begin
              dma2mem[49][25].run()  ;
            end

            begin
              gen[49][26].run()  ;
            end
            begin
              drv[49][26].run()  ;
            end
            begin
              dma2mem[49][26].run()  ;
            end

            begin
              gen[49][27].run()  ;
            end
            begin
              drv[49][27].run()  ;
            end
            begin
              dma2mem[49][27].run()  ;
            end

            begin
              gen[49][28].run()  ;
            end
            begin
              drv[49][28].run()  ;
            end
            begin
              dma2mem[49][28].run()  ;
            end

            begin
              gen[49][29].run()  ;
            end
            begin
              drv[49][29].run()  ;
            end
            begin
              dma2mem[49][29].run()  ;
            end

            begin
              gen[49][30].run()  ;
            end
            begin
              drv[49][30].run()  ;
            end
            begin
              dma2mem[49][30].run()  ;
            end

            begin
              gen[49][31].run()  ;
            end
            begin
              drv[49][31].run()  ;
            end
            begin
              dma2mem[49][31].run()  ;
            end

            begin
              gen[50][0].run()  ;
            end
            begin
              drv[50][0].run()  ;
            end
            begin
              dma2mem[50][0].run()  ;
            end

            begin
              gen[50][1].run()  ;
            end
            begin
              drv[50][1].run()  ;
            end
            begin
              dma2mem[50][1].run()  ;
            end

            begin
              gen[50][2].run()  ;
            end
            begin
              drv[50][2].run()  ;
            end
            begin
              dma2mem[50][2].run()  ;
            end

            begin
              gen[50][3].run()  ;
            end
            begin
              drv[50][3].run()  ;
            end
            begin
              dma2mem[50][3].run()  ;
            end

            begin
              gen[50][4].run()  ;
            end
            begin
              drv[50][4].run()  ;
            end
            begin
              dma2mem[50][4].run()  ;
            end

            begin
              gen[50][5].run()  ;
            end
            begin
              drv[50][5].run()  ;
            end
            begin
              dma2mem[50][5].run()  ;
            end

            begin
              gen[50][6].run()  ;
            end
            begin
              drv[50][6].run()  ;
            end
            begin
              dma2mem[50][6].run()  ;
            end

            begin
              gen[50][7].run()  ;
            end
            begin
              drv[50][7].run()  ;
            end
            begin
              dma2mem[50][7].run()  ;
            end

            begin
              gen[50][8].run()  ;
            end
            begin
              drv[50][8].run()  ;
            end
            begin
              dma2mem[50][8].run()  ;
            end

            begin
              gen[50][9].run()  ;
            end
            begin
              drv[50][9].run()  ;
            end
            begin
              dma2mem[50][9].run()  ;
            end

            begin
              gen[50][10].run()  ;
            end
            begin
              drv[50][10].run()  ;
            end
            begin
              dma2mem[50][10].run()  ;
            end

            begin
              gen[50][11].run()  ;
            end
            begin
              drv[50][11].run()  ;
            end
            begin
              dma2mem[50][11].run()  ;
            end

            begin
              gen[50][12].run()  ;
            end
            begin
              drv[50][12].run()  ;
            end
            begin
              dma2mem[50][12].run()  ;
            end

            begin
              gen[50][13].run()  ;
            end
            begin
              drv[50][13].run()  ;
            end
            begin
              dma2mem[50][13].run()  ;
            end

            begin
              gen[50][14].run()  ;
            end
            begin
              drv[50][14].run()  ;
            end
            begin
              dma2mem[50][14].run()  ;
            end

            begin
              gen[50][15].run()  ;
            end
            begin
              drv[50][15].run()  ;
            end
            begin
              dma2mem[50][15].run()  ;
            end

            begin
              gen[50][16].run()  ;
            end
            begin
              drv[50][16].run()  ;
            end
            begin
              dma2mem[50][16].run()  ;
            end

            begin
              gen[50][17].run()  ;
            end
            begin
              drv[50][17].run()  ;
            end
            begin
              dma2mem[50][17].run()  ;
            end

            begin
              gen[50][18].run()  ;
            end
            begin
              drv[50][18].run()  ;
            end
            begin
              dma2mem[50][18].run()  ;
            end

            begin
              gen[50][19].run()  ;
            end
            begin
              drv[50][19].run()  ;
            end
            begin
              dma2mem[50][19].run()  ;
            end

            begin
              gen[50][20].run()  ;
            end
            begin
              drv[50][20].run()  ;
            end
            begin
              dma2mem[50][20].run()  ;
            end

            begin
              gen[50][21].run()  ;
            end
            begin
              drv[50][21].run()  ;
            end
            begin
              dma2mem[50][21].run()  ;
            end

            begin
              gen[50][22].run()  ;
            end
            begin
              drv[50][22].run()  ;
            end
            begin
              dma2mem[50][22].run()  ;
            end

            begin
              gen[50][23].run()  ;
            end
            begin
              drv[50][23].run()  ;
            end
            begin
              dma2mem[50][23].run()  ;
            end

            begin
              gen[50][24].run()  ;
            end
            begin
              drv[50][24].run()  ;
            end
            begin
              dma2mem[50][24].run()  ;
            end

            begin
              gen[50][25].run()  ;
            end
            begin
              drv[50][25].run()  ;
            end
            begin
              dma2mem[50][25].run()  ;
            end

            begin
              gen[50][26].run()  ;
            end
            begin
              drv[50][26].run()  ;
            end
            begin
              dma2mem[50][26].run()  ;
            end

            begin
              gen[50][27].run()  ;
            end
            begin
              drv[50][27].run()  ;
            end
            begin
              dma2mem[50][27].run()  ;
            end

            begin
              gen[50][28].run()  ;
            end
            begin
              drv[50][28].run()  ;
            end
            begin
              dma2mem[50][28].run()  ;
            end

            begin
              gen[50][29].run()  ;
            end
            begin
              drv[50][29].run()  ;
            end
            begin
              dma2mem[50][29].run()  ;
            end

            begin
              gen[50][30].run()  ;
            end
            begin
              drv[50][30].run()  ;
            end
            begin
              dma2mem[50][30].run()  ;
            end

            begin
              gen[50][31].run()  ;
            end
            begin
              drv[50][31].run()  ;
            end
            begin
              dma2mem[50][31].run()  ;
            end

            begin
              gen[51][0].run()  ;
            end
            begin
              drv[51][0].run()  ;
            end
            begin
              dma2mem[51][0].run()  ;
            end

            begin
              gen[51][1].run()  ;
            end
            begin
              drv[51][1].run()  ;
            end
            begin
              dma2mem[51][1].run()  ;
            end

            begin
              gen[51][2].run()  ;
            end
            begin
              drv[51][2].run()  ;
            end
            begin
              dma2mem[51][2].run()  ;
            end

            begin
              gen[51][3].run()  ;
            end
            begin
              drv[51][3].run()  ;
            end
            begin
              dma2mem[51][3].run()  ;
            end

            begin
              gen[51][4].run()  ;
            end
            begin
              drv[51][4].run()  ;
            end
            begin
              dma2mem[51][4].run()  ;
            end

            begin
              gen[51][5].run()  ;
            end
            begin
              drv[51][5].run()  ;
            end
            begin
              dma2mem[51][5].run()  ;
            end

            begin
              gen[51][6].run()  ;
            end
            begin
              drv[51][6].run()  ;
            end
            begin
              dma2mem[51][6].run()  ;
            end

            begin
              gen[51][7].run()  ;
            end
            begin
              drv[51][7].run()  ;
            end
            begin
              dma2mem[51][7].run()  ;
            end

            begin
              gen[51][8].run()  ;
            end
            begin
              drv[51][8].run()  ;
            end
            begin
              dma2mem[51][8].run()  ;
            end

            begin
              gen[51][9].run()  ;
            end
            begin
              drv[51][9].run()  ;
            end
            begin
              dma2mem[51][9].run()  ;
            end

            begin
              gen[51][10].run()  ;
            end
            begin
              drv[51][10].run()  ;
            end
            begin
              dma2mem[51][10].run()  ;
            end

            begin
              gen[51][11].run()  ;
            end
            begin
              drv[51][11].run()  ;
            end
            begin
              dma2mem[51][11].run()  ;
            end

            begin
              gen[51][12].run()  ;
            end
            begin
              drv[51][12].run()  ;
            end
            begin
              dma2mem[51][12].run()  ;
            end

            begin
              gen[51][13].run()  ;
            end
            begin
              drv[51][13].run()  ;
            end
            begin
              dma2mem[51][13].run()  ;
            end

            begin
              gen[51][14].run()  ;
            end
            begin
              drv[51][14].run()  ;
            end
            begin
              dma2mem[51][14].run()  ;
            end

            begin
              gen[51][15].run()  ;
            end
            begin
              drv[51][15].run()  ;
            end
            begin
              dma2mem[51][15].run()  ;
            end

            begin
              gen[51][16].run()  ;
            end
            begin
              drv[51][16].run()  ;
            end
            begin
              dma2mem[51][16].run()  ;
            end

            begin
              gen[51][17].run()  ;
            end
            begin
              drv[51][17].run()  ;
            end
            begin
              dma2mem[51][17].run()  ;
            end

            begin
              gen[51][18].run()  ;
            end
            begin
              drv[51][18].run()  ;
            end
            begin
              dma2mem[51][18].run()  ;
            end

            begin
              gen[51][19].run()  ;
            end
            begin
              drv[51][19].run()  ;
            end
            begin
              dma2mem[51][19].run()  ;
            end

            begin
              gen[51][20].run()  ;
            end
            begin
              drv[51][20].run()  ;
            end
            begin
              dma2mem[51][20].run()  ;
            end

            begin
              gen[51][21].run()  ;
            end
            begin
              drv[51][21].run()  ;
            end
            begin
              dma2mem[51][21].run()  ;
            end

            begin
              gen[51][22].run()  ;
            end
            begin
              drv[51][22].run()  ;
            end
            begin
              dma2mem[51][22].run()  ;
            end

            begin
              gen[51][23].run()  ;
            end
            begin
              drv[51][23].run()  ;
            end
            begin
              dma2mem[51][23].run()  ;
            end

            begin
              gen[51][24].run()  ;
            end
            begin
              drv[51][24].run()  ;
            end
            begin
              dma2mem[51][24].run()  ;
            end

            begin
              gen[51][25].run()  ;
            end
            begin
              drv[51][25].run()  ;
            end
            begin
              dma2mem[51][25].run()  ;
            end

            begin
              gen[51][26].run()  ;
            end
            begin
              drv[51][26].run()  ;
            end
            begin
              dma2mem[51][26].run()  ;
            end

            begin
              gen[51][27].run()  ;
            end
            begin
              drv[51][27].run()  ;
            end
            begin
              dma2mem[51][27].run()  ;
            end

            begin
              gen[51][28].run()  ;
            end
            begin
              drv[51][28].run()  ;
            end
            begin
              dma2mem[51][28].run()  ;
            end

            begin
              gen[51][29].run()  ;
            end
            begin
              drv[51][29].run()  ;
            end
            begin
              dma2mem[51][29].run()  ;
            end

            begin
              gen[51][30].run()  ;
            end
            begin
              drv[51][30].run()  ;
            end
            begin
              dma2mem[51][30].run()  ;
            end

            begin
              gen[51][31].run()  ;
            end
            begin
              drv[51][31].run()  ;
            end
            begin
              dma2mem[51][31].run()  ;
            end

            begin
              gen[52][0].run()  ;
            end
            begin
              drv[52][0].run()  ;
            end
            begin
              dma2mem[52][0].run()  ;
            end

            begin
              gen[52][1].run()  ;
            end
            begin
              drv[52][1].run()  ;
            end
            begin
              dma2mem[52][1].run()  ;
            end

            begin
              gen[52][2].run()  ;
            end
            begin
              drv[52][2].run()  ;
            end
            begin
              dma2mem[52][2].run()  ;
            end

            begin
              gen[52][3].run()  ;
            end
            begin
              drv[52][3].run()  ;
            end
            begin
              dma2mem[52][3].run()  ;
            end

            begin
              gen[52][4].run()  ;
            end
            begin
              drv[52][4].run()  ;
            end
            begin
              dma2mem[52][4].run()  ;
            end

            begin
              gen[52][5].run()  ;
            end
            begin
              drv[52][5].run()  ;
            end
            begin
              dma2mem[52][5].run()  ;
            end

            begin
              gen[52][6].run()  ;
            end
            begin
              drv[52][6].run()  ;
            end
            begin
              dma2mem[52][6].run()  ;
            end

            begin
              gen[52][7].run()  ;
            end
            begin
              drv[52][7].run()  ;
            end
            begin
              dma2mem[52][7].run()  ;
            end

            begin
              gen[52][8].run()  ;
            end
            begin
              drv[52][8].run()  ;
            end
            begin
              dma2mem[52][8].run()  ;
            end

            begin
              gen[52][9].run()  ;
            end
            begin
              drv[52][9].run()  ;
            end
            begin
              dma2mem[52][9].run()  ;
            end

            begin
              gen[52][10].run()  ;
            end
            begin
              drv[52][10].run()  ;
            end
            begin
              dma2mem[52][10].run()  ;
            end

            begin
              gen[52][11].run()  ;
            end
            begin
              drv[52][11].run()  ;
            end
            begin
              dma2mem[52][11].run()  ;
            end

            begin
              gen[52][12].run()  ;
            end
            begin
              drv[52][12].run()  ;
            end
            begin
              dma2mem[52][12].run()  ;
            end

            begin
              gen[52][13].run()  ;
            end
            begin
              drv[52][13].run()  ;
            end
            begin
              dma2mem[52][13].run()  ;
            end

            begin
              gen[52][14].run()  ;
            end
            begin
              drv[52][14].run()  ;
            end
            begin
              dma2mem[52][14].run()  ;
            end

            begin
              gen[52][15].run()  ;
            end
            begin
              drv[52][15].run()  ;
            end
            begin
              dma2mem[52][15].run()  ;
            end

            begin
              gen[52][16].run()  ;
            end
            begin
              drv[52][16].run()  ;
            end
            begin
              dma2mem[52][16].run()  ;
            end

            begin
              gen[52][17].run()  ;
            end
            begin
              drv[52][17].run()  ;
            end
            begin
              dma2mem[52][17].run()  ;
            end

            begin
              gen[52][18].run()  ;
            end
            begin
              drv[52][18].run()  ;
            end
            begin
              dma2mem[52][18].run()  ;
            end

            begin
              gen[52][19].run()  ;
            end
            begin
              drv[52][19].run()  ;
            end
            begin
              dma2mem[52][19].run()  ;
            end

            begin
              gen[52][20].run()  ;
            end
            begin
              drv[52][20].run()  ;
            end
            begin
              dma2mem[52][20].run()  ;
            end

            begin
              gen[52][21].run()  ;
            end
            begin
              drv[52][21].run()  ;
            end
            begin
              dma2mem[52][21].run()  ;
            end

            begin
              gen[52][22].run()  ;
            end
            begin
              drv[52][22].run()  ;
            end
            begin
              dma2mem[52][22].run()  ;
            end

            begin
              gen[52][23].run()  ;
            end
            begin
              drv[52][23].run()  ;
            end
            begin
              dma2mem[52][23].run()  ;
            end

            begin
              gen[52][24].run()  ;
            end
            begin
              drv[52][24].run()  ;
            end
            begin
              dma2mem[52][24].run()  ;
            end

            begin
              gen[52][25].run()  ;
            end
            begin
              drv[52][25].run()  ;
            end
            begin
              dma2mem[52][25].run()  ;
            end

            begin
              gen[52][26].run()  ;
            end
            begin
              drv[52][26].run()  ;
            end
            begin
              dma2mem[52][26].run()  ;
            end

            begin
              gen[52][27].run()  ;
            end
            begin
              drv[52][27].run()  ;
            end
            begin
              dma2mem[52][27].run()  ;
            end

            begin
              gen[52][28].run()  ;
            end
            begin
              drv[52][28].run()  ;
            end
            begin
              dma2mem[52][28].run()  ;
            end

            begin
              gen[52][29].run()  ;
            end
            begin
              drv[52][29].run()  ;
            end
            begin
              dma2mem[52][29].run()  ;
            end

            begin
              gen[52][30].run()  ;
            end
            begin
              drv[52][30].run()  ;
            end
            begin
              dma2mem[52][30].run()  ;
            end

            begin
              gen[52][31].run()  ;
            end
            begin
              drv[52][31].run()  ;
            end
            begin
              dma2mem[52][31].run()  ;
            end

            begin
              gen[53][0].run()  ;
            end
            begin
              drv[53][0].run()  ;
            end
            begin
              dma2mem[53][0].run()  ;
            end

            begin
              gen[53][1].run()  ;
            end
            begin
              drv[53][1].run()  ;
            end
            begin
              dma2mem[53][1].run()  ;
            end

            begin
              gen[53][2].run()  ;
            end
            begin
              drv[53][2].run()  ;
            end
            begin
              dma2mem[53][2].run()  ;
            end

            begin
              gen[53][3].run()  ;
            end
            begin
              drv[53][3].run()  ;
            end
            begin
              dma2mem[53][3].run()  ;
            end

            begin
              gen[53][4].run()  ;
            end
            begin
              drv[53][4].run()  ;
            end
            begin
              dma2mem[53][4].run()  ;
            end

            begin
              gen[53][5].run()  ;
            end
            begin
              drv[53][5].run()  ;
            end
            begin
              dma2mem[53][5].run()  ;
            end

            begin
              gen[53][6].run()  ;
            end
            begin
              drv[53][6].run()  ;
            end
            begin
              dma2mem[53][6].run()  ;
            end

            begin
              gen[53][7].run()  ;
            end
            begin
              drv[53][7].run()  ;
            end
            begin
              dma2mem[53][7].run()  ;
            end

            begin
              gen[53][8].run()  ;
            end
            begin
              drv[53][8].run()  ;
            end
            begin
              dma2mem[53][8].run()  ;
            end

            begin
              gen[53][9].run()  ;
            end
            begin
              drv[53][9].run()  ;
            end
            begin
              dma2mem[53][9].run()  ;
            end

            begin
              gen[53][10].run()  ;
            end
            begin
              drv[53][10].run()  ;
            end
            begin
              dma2mem[53][10].run()  ;
            end

            begin
              gen[53][11].run()  ;
            end
            begin
              drv[53][11].run()  ;
            end
            begin
              dma2mem[53][11].run()  ;
            end

            begin
              gen[53][12].run()  ;
            end
            begin
              drv[53][12].run()  ;
            end
            begin
              dma2mem[53][12].run()  ;
            end

            begin
              gen[53][13].run()  ;
            end
            begin
              drv[53][13].run()  ;
            end
            begin
              dma2mem[53][13].run()  ;
            end

            begin
              gen[53][14].run()  ;
            end
            begin
              drv[53][14].run()  ;
            end
            begin
              dma2mem[53][14].run()  ;
            end

            begin
              gen[53][15].run()  ;
            end
            begin
              drv[53][15].run()  ;
            end
            begin
              dma2mem[53][15].run()  ;
            end

            begin
              gen[53][16].run()  ;
            end
            begin
              drv[53][16].run()  ;
            end
            begin
              dma2mem[53][16].run()  ;
            end

            begin
              gen[53][17].run()  ;
            end
            begin
              drv[53][17].run()  ;
            end
            begin
              dma2mem[53][17].run()  ;
            end

            begin
              gen[53][18].run()  ;
            end
            begin
              drv[53][18].run()  ;
            end
            begin
              dma2mem[53][18].run()  ;
            end

            begin
              gen[53][19].run()  ;
            end
            begin
              drv[53][19].run()  ;
            end
            begin
              dma2mem[53][19].run()  ;
            end

            begin
              gen[53][20].run()  ;
            end
            begin
              drv[53][20].run()  ;
            end
            begin
              dma2mem[53][20].run()  ;
            end

            begin
              gen[53][21].run()  ;
            end
            begin
              drv[53][21].run()  ;
            end
            begin
              dma2mem[53][21].run()  ;
            end

            begin
              gen[53][22].run()  ;
            end
            begin
              drv[53][22].run()  ;
            end
            begin
              dma2mem[53][22].run()  ;
            end

            begin
              gen[53][23].run()  ;
            end
            begin
              drv[53][23].run()  ;
            end
            begin
              dma2mem[53][23].run()  ;
            end

            begin
              gen[53][24].run()  ;
            end
            begin
              drv[53][24].run()  ;
            end
            begin
              dma2mem[53][24].run()  ;
            end

            begin
              gen[53][25].run()  ;
            end
            begin
              drv[53][25].run()  ;
            end
            begin
              dma2mem[53][25].run()  ;
            end

            begin
              gen[53][26].run()  ;
            end
            begin
              drv[53][26].run()  ;
            end
            begin
              dma2mem[53][26].run()  ;
            end

            begin
              gen[53][27].run()  ;
            end
            begin
              drv[53][27].run()  ;
            end
            begin
              dma2mem[53][27].run()  ;
            end

            begin
              gen[53][28].run()  ;
            end
            begin
              drv[53][28].run()  ;
            end
            begin
              dma2mem[53][28].run()  ;
            end

            begin
              gen[53][29].run()  ;
            end
            begin
              drv[53][29].run()  ;
            end
            begin
              dma2mem[53][29].run()  ;
            end

            begin
              gen[53][30].run()  ;
            end
            begin
              drv[53][30].run()  ;
            end
            begin
              dma2mem[53][30].run()  ;
            end

            begin
              gen[53][31].run()  ;
            end
            begin
              drv[53][31].run()  ;
            end
            begin
              dma2mem[53][31].run()  ;
            end

            begin
              gen[54][0].run()  ;
            end
            begin
              drv[54][0].run()  ;
            end
            begin
              dma2mem[54][0].run()  ;
            end

            begin
              gen[54][1].run()  ;
            end
            begin
              drv[54][1].run()  ;
            end
            begin
              dma2mem[54][1].run()  ;
            end

            begin
              gen[54][2].run()  ;
            end
            begin
              drv[54][2].run()  ;
            end
            begin
              dma2mem[54][2].run()  ;
            end

            begin
              gen[54][3].run()  ;
            end
            begin
              drv[54][3].run()  ;
            end
            begin
              dma2mem[54][3].run()  ;
            end

            begin
              gen[54][4].run()  ;
            end
            begin
              drv[54][4].run()  ;
            end
            begin
              dma2mem[54][4].run()  ;
            end

            begin
              gen[54][5].run()  ;
            end
            begin
              drv[54][5].run()  ;
            end
            begin
              dma2mem[54][5].run()  ;
            end

            begin
              gen[54][6].run()  ;
            end
            begin
              drv[54][6].run()  ;
            end
            begin
              dma2mem[54][6].run()  ;
            end

            begin
              gen[54][7].run()  ;
            end
            begin
              drv[54][7].run()  ;
            end
            begin
              dma2mem[54][7].run()  ;
            end

            begin
              gen[54][8].run()  ;
            end
            begin
              drv[54][8].run()  ;
            end
            begin
              dma2mem[54][8].run()  ;
            end

            begin
              gen[54][9].run()  ;
            end
            begin
              drv[54][9].run()  ;
            end
            begin
              dma2mem[54][9].run()  ;
            end

            begin
              gen[54][10].run()  ;
            end
            begin
              drv[54][10].run()  ;
            end
            begin
              dma2mem[54][10].run()  ;
            end

            begin
              gen[54][11].run()  ;
            end
            begin
              drv[54][11].run()  ;
            end
            begin
              dma2mem[54][11].run()  ;
            end

            begin
              gen[54][12].run()  ;
            end
            begin
              drv[54][12].run()  ;
            end
            begin
              dma2mem[54][12].run()  ;
            end

            begin
              gen[54][13].run()  ;
            end
            begin
              drv[54][13].run()  ;
            end
            begin
              dma2mem[54][13].run()  ;
            end

            begin
              gen[54][14].run()  ;
            end
            begin
              drv[54][14].run()  ;
            end
            begin
              dma2mem[54][14].run()  ;
            end

            begin
              gen[54][15].run()  ;
            end
            begin
              drv[54][15].run()  ;
            end
            begin
              dma2mem[54][15].run()  ;
            end

            begin
              gen[54][16].run()  ;
            end
            begin
              drv[54][16].run()  ;
            end
            begin
              dma2mem[54][16].run()  ;
            end

            begin
              gen[54][17].run()  ;
            end
            begin
              drv[54][17].run()  ;
            end
            begin
              dma2mem[54][17].run()  ;
            end

            begin
              gen[54][18].run()  ;
            end
            begin
              drv[54][18].run()  ;
            end
            begin
              dma2mem[54][18].run()  ;
            end

            begin
              gen[54][19].run()  ;
            end
            begin
              drv[54][19].run()  ;
            end
            begin
              dma2mem[54][19].run()  ;
            end

            begin
              gen[54][20].run()  ;
            end
            begin
              drv[54][20].run()  ;
            end
            begin
              dma2mem[54][20].run()  ;
            end

            begin
              gen[54][21].run()  ;
            end
            begin
              drv[54][21].run()  ;
            end
            begin
              dma2mem[54][21].run()  ;
            end

            begin
              gen[54][22].run()  ;
            end
            begin
              drv[54][22].run()  ;
            end
            begin
              dma2mem[54][22].run()  ;
            end

            begin
              gen[54][23].run()  ;
            end
            begin
              drv[54][23].run()  ;
            end
            begin
              dma2mem[54][23].run()  ;
            end

            begin
              gen[54][24].run()  ;
            end
            begin
              drv[54][24].run()  ;
            end
            begin
              dma2mem[54][24].run()  ;
            end

            begin
              gen[54][25].run()  ;
            end
            begin
              drv[54][25].run()  ;
            end
            begin
              dma2mem[54][25].run()  ;
            end

            begin
              gen[54][26].run()  ;
            end
            begin
              drv[54][26].run()  ;
            end
            begin
              dma2mem[54][26].run()  ;
            end

            begin
              gen[54][27].run()  ;
            end
            begin
              drv[54][27].run()  ;
            end
            begin
              dma2mem[54][27].run()  ;
            end

            begin
              gen[54][28].run()  ;
            end
            begin
              drv[54][28].run()  ;
            end
            begin
              dma2mem[54][28].run()  ;
            end

            begin
              gen[54][29].run()  ;
            end
            begin
              drv[54][29].run()  ;
            end
            begin
              dma2mem[54][29].run()  ;
            end

            begin
              gen[54][30].run()  ;
            end
            begin
              drv[54][30].run()  ;
            end
            begin
              dma2mem[54][30].run()  ;
            end

            begin
              gen[54][31].run()  ;
            end
            begin
              drv[54][31].run()  ;
            end
            begin
              dma2mem[54][31].run()  ;
            end

            begin
              gen[55][0].run()  ;
            end
            begin
              drv[55][0].run()  ;
            end
            begin
              dma2mem[55][0].run()  ;
            end

            begin
              gen[55][1].run()  ;
            end
            begin
              drv[55][1].run()  ;
            end
            begin
              dma2mem[55][1].run()  ;
            end

            begin
              gen[55][2].run()  ;
            end
            begin
              drv[55][2].run()  ;
            end
            begin
              dma2mem[55][2].run()  ;
            end

            begin
              gen[55][3].run()  ;
            end
            begin
              drv[55][3].run()  ;
            end
            begin
              dma2mem[55][3].run()  ;
            end

            begin
              gen[55][4].run()  ;
            end
            begin
              drv[55][4].run()  ;
            end
            begin
              dma2mem[55][4].run()  ;
            end

            begin
              gen[55][5].run()  ;
            end
            begin
              drv[55][5].run()  ;
            end
            begin
              dma2mem[55][5].run()  ;
            end

            begin
              gen[55][6].run()  ;
            end
            begin
              drv[55][6].run()  ;
            end
            begin
              dma2mem[55][6].run()  ;
            end

            begin
              gen[55][7].run()  ;
            end
            begin
              drv[55][7].run()  ;
            end
            begin
              dma2mem[55][7].run()  ;
            end

            begin
              gen[55][8].run()  ;
            end
            begin
              drv[55][8].run()  ;
            end
            begin
              dma2mem[55][8].run()  ;
            end

            begin
              gen[55][9].run()  ;
            end
            begin
              drv[55][9].run()  ;
            end
            begin
              dma2mem[55][9].run()  ;
            end

            begin
              gen[55][10].run()  ;
            end
            begin
              drv[55][10].run()  ;
            end
            begin
              dma2mem[55][10].run()  ;
            end

            begin
              gen[55][11].run()  ;
            end
            begin
              drv[55][11].run()  ;
            end
            begin
              dma2mem[55][11].run()  ;
            end

            begin
              gen[55][12].run()  ;
            end
            begin
              drv[55][12].run()  ;
            end
            begin
              dma2mem[55][12].run()  ;
            end

            begin
              gen[55][13].run()  ;
            end
            begin
              drv[55][13].run()  ;
            end
            begin
              dma2mem[55][13].run()  ;
            end

            begin
              gen[55][14].run()  ;
            end
            begin
              drv[55][14].run()  ;
            end
            begin
              dma2mem[55][14].run()  ;
            end

            begin
              gen[55][15].run()  ;
            end
            begin
              drv[55][15].run()  ;
            end
            begin
              dma2mem[55][15].run()  ;
            end

            begin
              gen[55][16].run()  ;
            end
            begin
              drv[55][16].run()  ;
            end
            begin
              dma2mem[55][16].run()  ;
            end

            begin
              gen[55][17].run()  ;
            end
            begin
              drv[55][17].run()  ;
            end
            begin
              dma2mem[55][17].run()  ;
            end

            begin
              gen[55][18].run()  ;
            end
            begin
              drv[55][18].run()  ;
            end
            begin
              dma2mem[55][18].run()  ;
            end

            begin
              gen[55][19].run()  ;
            end
            begin
              drv[55][19].run()  ;
            end
            begin
              dma2mem[55][19].run()  ;
            end

            begin
              gen[55][20].run()  ;
            end
            begin
              drv[55][20].run()  ;
            end
            begin
              dma2mem[55][20].run()  ;
            end

            begin
              gen[55][21].run()  ;
            end
            begin
              drv[55][21].run()  ;
            end
            begin
              dma2mem[55][21].run()  ;
            end

            begin
              gen[55][22].run()  ;
            end
            begin
              drv[55][22].run()  ;
            end
            begin
              dma2mem[55][22].run()  ;
            end

            begin
              gen[55][23].run()  ;
            end
            begin
              drv[55][23].run()  ;
            end
            begin
              dma2mem[55][23].run()  ;
            end

            begin
              gen[55][24].run()  ;
            end
            begin
              drv[55][24].run()  ;
            end
            begin
              dma2mem[55][24].run()  ;
            end

            begin
              gen[55][25].run()  ;
            end
            begin
              drv[55][25].run()  ;
            end
            begin
              dma2mem[55][25].run()  ;
            end

            begin
              gen[55][26].run()  ;
            end
            begin
              drv[55][26].run()  ;
            end
            begin
              dma2mem[55][26].run()  ;
            end

            begin
              gen[55][27].run()  ;
            end
            begin
              drv[55][27].run()  ;
            end
            begin
              dma2mem[55][27].run()  ;
            end

            begin
              gen[55][28].run()  ;
            end
            begin
              drv[55][28].run()  ;
            end
            begin
              dma2mem[55][28].run()  ;
            end

            begin
              gen[55][29].run()  ;
            end
            begin
              drv[55][29].run()  ;
            end
            begin
              dma2mem[55][29].run()  ;
            end

            begin
              gen[55][30].run()  ;
            end
            begin
              drv[55][30].run()  ;
            end
            begin
              dma2mem[55][30].run()  ;
            end

            begin
              gen[55][31].run()  ;
            end
            begin
              drv[55][31].run()  ;
            end
            begin
              dma2mem[55][31].run()  ;
            end

            begin
              gen[56][0].run()  ;
            end
            begin
              drv[56][0].run()  ;
            end
            begin
              dma2mem[56][0].run()  ;
            end

            begin
              gen[56][1].run()  ;
            end
            begin
              drv[56][1].run()  ;
            end
            begin
              dma2mem[56][1].run()  ;
            end

            begin
              gen[56][2].run()  ;
            end
            begin
              drv[56][2].run()  ;
            end
            begin
              dma2mem[56][2].run()  ;
            end

            begin
              gen[56][3].run()  ;
            end
            begin
              drv[56][3].run()  ;
            end
            begin
              dma2mem[56][3].run()  ;
            end

            begin
              gen[56][4].run()  ;
            end
            begin
              drv[56][4].run()  ;
            end
            begin
              dma2mem[56][4].run()  ;
            end

            begin
              gen[56][5].run()  ;
            end
            begin
              drv[56][5].run()  ;
            end
            begin
              dma2mem[56][5].run()  ;
            end

            begin
              gen[56][6].run()  ;
            end
            begin
              drv[56][6].run()  ;
            end
            begin
              dma2mem[56][6].run()  ;
            end

            begin
              gen[56][7].run()  ;
            end
            begin
              drv[56][7].run()  ;
            end
            begin
              dma2mem[56][7].run()  ;
            end

            begin
              gen[56][8].run()  ;
            end
            begin
              drv[56][8].run()  ;
            end
            begin
              dma2mem[56][8].run()  ;
            end

            begin
              gen[56][9].run()  ;
            end
            begin
              drv[56][9].run()  ;
            end
            begin
              dma2mem[56][9].run()  ;
            end

            begin
              gen[56][10].run()  ;
            end
            begin
              drv[56][10].run()  ;
            end
            begin
              dma2mem[56][10].run()  ;
            end

            begin
              gen[56][11].run()  ;
            end
            begin
              drv[56][11].run()  ;
            end
            begin
              dma2mem[56][11].run()  ;
            end

            begin
              gen[56][12].run()  ;
            end
            begin
              drv[56][12].run()  ;
            end
            begin
              dma2mem[56][12].run()  ;
            end

            begin
              gen[56][13].run()  ;
            end
            begin
              drv[56][13].run()  ;
            end
            begin
              dma2mem[56][13].run()  ;
            end

            begin
              gen[56][14].run()  ;
            end
            begin
              drv[56][14].run()  ;
            end
            begin
              dma2mem[56][14].run()  ;
            end

            begin
              gen[56][15].run()  ;
            end
            begin
              drv[56][15].run()  ;
            end
            begin
              dma2mem[56][15].run()  ;
            end

            begin
              gen[56][16].run()  ;
            end
            begin
              drv[56][16].run()  ;
            end
            begin
              dma2mem[56][16].run()  ;
            end

            begin
              gen[56][17].run()  ;
            end
            begin
              drv[56][17].run()  ;
            end
            begin
              dma2mem[56][17].run()  ;
            end

            begin
              gen[56][18].run()  ;
            end
            begin
              drv[56][18].run()  ;
            end
            begin
              dma2mem[56][18].run()  ;
            end

            begin
              gen[56][19].run()  ;
            end
            begin
              drv[56][19].run()  ;
            end
            begin
              dma2mem[56][19].run()  ;
            end

            begin
              gen[56][20].run()  ;
            end
            begin
              drv[56][20].run()  ;
            end
            begin
              dma2mem[56][20].run()  ;
            end

            begin
              gen[56][21].run()  ;
            end
            begin
              drv[56][21].run()  ;
            end
            begin
              dma2mem[56][21].run()  ;
            end

            begin
              gen[56][22].run()  ;
            end
            begin
              drv[56][22].run()  ;
            end
            begin
              dma2mem[56][22].run()  ;
            end

            begin
              gen[56][23].run()  ;
            end
            begin
              drv[56][23].run()  ;
            end
            begin
              dma2mem[56][23].run()  ;
            end

            begin
              gen[56][24].run()  ;
            end
            begin
              drv[56][24].run()  ;
            end
            begin
              dma2mem[56][24].run()  ;
            end

            begin
              gen[56][25].run()  ;
            end
            begin
              drv[56][25].run()  ;
            end
            begin
              dma2mem[56][25].run()  ;
            end

            begin
              gen[56][26].run()  ;
            end
            begin
              drv[56][26].run()  ;
            end
            begin
              dma2mem[56][26].run()  ;
            end

            begin
              gen[56][27].run()  ;
            end
            begin
              drv[56][27].run()  ;
            end
            begin
              dma2mem[56][27].run()  ;
            end

            begin
              gen[56][28].run()  ;
            end
            begin
              drv[56][28].run()  ;
            end
            begin
              dma2mem[56][28].run()  ;
            end

            begin
              gen[56][29].run()  ;
            end
            begin
              drv[56][29].run()  ;
            end
            begin
              dma2mem[56][29].run()  ;
            end

            begin
              gen[56][30].run()  ;
            end
            begin
              drv[56][30].run()  ;
            end
            begin
              dma2mem[56][30].run()  ;
            end

            begin
              gen[56][31].run()  ;
            end
            begin
              drv[56][31].run()  ;
            end
            begin
              dma2mem[56][31].run()  ;
            end

            begin
              gen[57][0].run()  ;
            end
            begin
              drv[57][0].run()  ;
            end
            begin
              dma2mem[57][0].run()  ;
            end

            begin
              gen[57][1].run()  ;
            end
            begin
              drv[57][1].run()  ;
            end
            begin
              dma2mem[57][1].run()  ;
            end

            begin
              gen[57][2].run()  ;
            end
            begin
              drv[57][2].run()  ;
            end
            begin
              dma2mem[57][2].run()  ;
            end

            begin
              gen[57][3].run()  ;
            end
            begin
              drv[57][3].run()  ;
            end
            begin
              dma2mem[57][3].run()  ;
            end

            begin
              gen[57][4].run()  ;
            end
            begin
              drv[57][4].run()  ;
            end
            begin
              dma2mem[57][4].run()  ;
            end

            begin
              gen[57][5].run()  ;
            end
            begin
              drv[57][5].run()  ;
            end
            begin
              dma2mem[57][5].run()  ;
            end

            begin
              gen[57][6].run()  ;
            end
            begin
              drv[57][6].run()  ;
            end
            begin
              dma2mem[57][6].run()  ;
            end

            begin
              gen[57][7].run()  ;
            end
            begin
              drv[57][7].run()  ;
            end
            begin
              dma2mem[57][7].run()  ;
            end

            begin
              gen[57][8].run()  ;
            end
            begin
              drv[57][8].run()  ;
            end
            begin
              dma2mem[57][8].run()  ;
            end

            begin
              gen[57][9].run()  ;
            end
            begin
              drv[57][9].run()  ;
            end
            begin
              dma2mem[57][9].run()  ;
            end

            begin
              gen[57][10].run()  ;
            end
            begin
              drv[57][10].run()  ;
            end
            begin
              dma2mem[57][10].run()  ;
            end

            begin
              gen[57][11].run()  ;
            end
            begin
              drv[57][11].run()  ;
            end
            begin
              dma2mem[57][11].run()  ;
            end

            begin
              gen[57][12].run()  ;
            end
            begin
              drv[57][12].run()  ;
            end
            begin
              dma2mem[57][12].run()  ;
            end

            begin
              gen[57][13].run()  ;
            end
            begin
              drv[57][13].run()  ;
            end
            begin
              dma2mem[57][13].run()  ;
            end

            begin
              gen[57][14].run()  ;
            end
            begin
              drv[57][14].run()  ;
            end
            begin
              dma2mem[57][14].run()  ;
            end

            begin
              gen[57][15].run()  ;
            end
            begin
              drv[57][15].run()  ;
            end
            begin
              dma2mem[57][15].run()  ;
            end

            begin
              gen[57][16].run()  ;
            end
            begin
              drv[57][16].run()  ;
            end
            begin
              dma2mem[57][16].run()  ;
            end

            begin
              gen[57][17].run()  ;
            end
            begin
              drv[57][17].run()  ;
            end
            begin
              dma2mem[57][17].run()  ;
            end

            begin
              gen[57][18].run()  ;
            end
            begin
              drv[57][18].run()  ;
            end
            begin
              dma2mem[57][18].run()  ;
            end

            begin
              gen[57][19].run()  ;
            end
            begin
              drv[57][19].run()  ;
            end
            begin
              dma2mem[57][19].run()  ;
            end

            begin
              gen[57][20].run()  ;
            end
            begin
              drv[57][20].run()  ;
            end
            begin
              dma2mem[57][20].run()  ;
            end

            begin
              gen[57][21].run()  ;
            end
            begin
              drv[57][21].run()  ;
            end
            begin
              dma2mem[57][21].run()  ;
            end

            begin
              gen[57][22].run()  ;
            end
            begin
              drv[57][22].run()  ;
            end
            begin
              dma2mem[57][22].run()  ;
            end

            begin
              gen[57][23].run()  ;
            end
            begin
              drv[57][23].run()  ;
            end
            begin
              dma2mem[57][23].run()  ;
            end

            begin
              gen[57][24].run()  ;
            end
            begin
              drv[57][24].run()  ;
            end
            begin
              dma2mem[57][24].run()  ;
            end

            begin
              gen[57][25].run()  ;
            end
            begin
              drv[57][25].run()  ;
            end
            begin
              dma2mem[57][25].run()  ;
            end

            begin
              gen[57][26].run()  ;
            end
            begin
              drv[57][26].run()  ;
            end
            begin
              dma2mem[57][26].run()  ;
            end

            begin
              gen[57][27].run()  ;
            end
            begin
              drv[57][27].run()  ;
            end
            begin
              dma2mem[57][27].run()  ;
            end

            begin
              gen[57][28].run()  ;
            end
            begin
              drv[57][28].run()  ;
            end
            begin
              dma2mem[57][28].run()  ;
            end

            begin
              gen[57][29].run()  ;
            end
            begin
              drv[57][29].run()  ;
            end
            begin
              dma2mem[57][29].run()  ;
            end

            begin
              gen[57][30].run()  ;
            end
            begin
              drv[57][30].run()  ;
            end
            begin
              dma2mem[57][30].run()  ;
            end

            begin
              gen[57][31].run()  ;
            end
            begin
              drv[57][31].run()  ;
            end
            begin
              dma2mem[57][31].run()  ;
            end

            begin
              gen[58][0].run()  ;
            end
            begin
              drv[58][0].run()  ;
            end
            begin
              dma2mem[58][0].run()  ;
            end

            begin
              gen[58][1].run()  ;
            end
            begin
              drv[58][1].run()  ;
            end
            begin
              dma2mem[58][1].run()  ;
            end

            begin
              gen[58][2].run()  ;
            end
            begin
              drv[58][2].run()  ;
            end
            begin
              dma2mem[58][2].run()  ;
            end

            begin
              gen[58][3].run()  ;
            end
            begin
              drv[58][3].run()  ;
            end
            begin
              dma2mem[58][3].run()  ;
            end

            begin
              gen[58][4].run()  ;
            end
            begin
              drv[58][4].run()  ;
            end
            begin
              dma2mem[58][4].run()  ;
            end

            begin
              gen[58][5].run()  ;
            end
            begin
              drv[58][5].run()  ;
            end
            begin
              dma2mem[58][5].run()  ;
            end

            begin
              gen[58][6].run()  ;
            end
            begin
              drv[58][6].run()  ;
            end
            begin
              dma2mem[58][6].run()  ;
            end

            begin
              gen[58][7].run()  ;
            end
            begin
              drv[58][7].run()  ;
            end
            begin
              dma2mem[58][7].run()  ;
            end

            begin
              gen[58][8].run()  ;
            end
            begin
              drv[58][8].run()  ;
            end
            begin
              dma2mem[58][8].run()  ;
            end

            begin
              gen[58][9].run()  ;
            end
            begin
              drv[58][9].run()  ;
            end
            begin
              dma2mem[58][9].run()  ;
            end

            begin
              gen[58][10].run()  ;
            end
            begin
              drv[58][10].run()  ;
            end
            begin
              dma2mem[58][10].run()  ;
            end

            begin
              gen[58][11].run()  ;
            end
            begin
              drv[58][11].run()  ;
            end
            begin
              dma2mem[58][11].run()  ;
            end

            begin
              gen[58][12].run()  ;
            end
            begin
              drv[58][12].run()  ;
            end
            begin
              dma2mem[58][12].run()  ;
            end

            begin
              gen[58][13].run()  ;
            end
            begin
              drv[58][13].run()  ;
            end
            begin
              dma2mem[58][13].run()  ;
            end

            begin
              gen[58][14].run()  ;
            end
            begin
              drv[58][14].run()  ;
            end
            begin
              dma2mem[58][14].run()  ;
            end

            begin
              gen[58][15].run()  ;
            end
            begin
              drv[58][15].run()  ;
            end
            begin
              dma2mem[58][15].run()  ;
            end

            begin
              gen[58][16].run()  ;
            end
            begin
              drv[58][16].run()  ;
            end
            begin
              dma2mem[58][16].run()  ;
            end

            begin
              gen[58][17].run()  ;
            end
            begin
              drv[58][17].run()  ;
            end
            begin
              dma2mem[58][17].run()  ;
            end

            begin
              gen[58][18].run()  ;
            end
            begin
              drv[58][18].run()  ;
            end
            begin
              dma2mem[58][18].run()  ;
            end

            begin
              gen[58][19].run()  ;
            end
            begin
              drv[58][19].run()  ;
            end
            begin
              dma2mem[58][19].run()  ;
            end

            begin
              gen[58][20].run()  ;
            end
            begin
              drv[58][20].run()  ;
            end
            begin
              dma2mem[58][20].run()  ;
            end

            begin
              gen[58][21].run()  ;
            end
            begin
              drv[58][21].run()  ;
            end
            begin
              dma2mem[58][21].run()  ;
            end

            begin
              gen[58][22].run()  ;
            end
            begin
              drv[58][22].run()  ;
            end
            begin
              dma2mem[58][22].run()  ;
            end

            begin
              gen[58][23].run()  ;
            end
            begin
              drv[58][23].run()  ;
            end
            begin
              dma2mem[58][23].run()  ;
            end

            begin
              gen[58][24].run()  ;
            end
            begin
              drv[58][24].run()  ;
            end
            begin
              dma2mem[58][24].run()  ;
            end

            begin
              gen[58][25].run()  ;
            end
            begin
              drv[58][25].run()  ;
            end
            begin
              dma2mem[58][25].run()  ;
            end

            begin
              gen[58][26].run()  ;
            end
            begin
              drv[58][26].run()  ;
            end
            begin
              dma2mem[58][26].run()  ;
            end

            begin
              gen[58][27].run()  ;
            end
            begin
              drv[58][27].run()  ;
            end
            begin
              dma2mem[58][27].run()  ;
            end

            begin
              gen[58][28].run()  ;
            end
            begin
              drv[58][28].run()  ;
            end
            begin
              dma2mem[58][28].run()  ;
            end

            begin
              gen[58][29].run()  ;
            end
            begin
              drv[58][29].run()  ;
            end
            begin
              dma2mem[58][29].run()  ;
            end

            begin
              gen[58][30].run()  ;
            end
            begin
              drv[58][30].run()  ;
            end
            begin
              dma2mem[58][30].run()  ;
            end

            begin
              gen[58][31].run()  ;
            end
            begin
              drv[58][31].run()  ;
            end
            begin
              dma2mem[58][31].run()  ;
            end

            begin
              gen[59][0].run()  ;
            end
            begin
              drv[59][0].run()  ;
            end
            begin
              dma2mem[59][0].run()  ;
            end

            begin
              gen[59][1].run()  ;
            end
            begin
              drv[59][1].run()  ;
            end
            begin
              dma2mem[59][1].run()  ;
            end

            begin
              gen[59][2].run()  ;
            end
            begin
              drv[59][2].run()  ;
            end
            begin
              dma2mem[59][2].run()  ;
            end

            begin
              gen[59][3].run()  ;
            end
            begin
              drv[59][3].run()  ;
            end
            begin
              dma2mem[59][3].run()  ;
            end

            begin
              gen[59][4].run()  ;
            end
            begin
              drv[59][4].run()  ;
            end
            begin
              dma2mem[59][4].run()  ;
            end

            begin
              gen[59][5].run()  ;
            end
            begin
              drv[59][5].run()  ;
            end
            begin
              dma2mem[59][5].run()  ;
            end

            begin
              gen[59][6].run()  ;
            end
            begin
              drv[59][6].run()  ;
            end
            begin
              dma2mem[59][6].run()  ;
            end

            begin
              gen[59][7].run()  ;
            end
            begin
              drv[59][7].run()  ;
            end
            begin
              dma2mem[59][7].run()  ;
            end

            begin
              gen[59][8].run()  ;
            end
            begin
              drv[59][8].run()  ;
            end
            begin
              dma2mem[59][8].run()  ;
            end

            begin
              gen[59][9].run()  ;
            end
            begin
              drv[59][9].run()  ;
            end
            begin
              dma2mem[59][9].run()  ;
            end

            begin
              gen[59][10].run()  ;
            end
            begin
              drv[59][10].run()  ;
            end
            begin
              dma2mem[59][10].run()  ;
            end

            begin
              gen[59][11].run()  ;
            end
            begin
              drv[59][11].run()  ;
            end
            begin
              dma2mem[59][11].run()  ;
            end

            begin
              gen[59][12].run()  ;
            end
            begin
              drv[59][12].run()  ;
            end
            begin
              dma2mem[59][12].run()  ;
            end

            begin
              gen[59][13].run()  ;
            end
            begin
              drv[59][13].run()  ;
            end
            begin
              dma2mem[59][13].run()  ;
            end

            begin
              gen[59][14].run()  ;
            end
            begin
              drv[59][14].run()  ;
            end
            begin
              dma2mem[59][14].run()  ;
            end

            begin
              gen[59][15].run()  ;
            end
            begin
              drv[59][15].run()  ;
            end
            begin
              dma2mem[59][15].run()  ;
            end

            begin
              gen[59][16].run()  ;
            end
            begin
              drv[59][16].run()  ;
            end
            begin
              dma2mem[59][16].run()  ;
            end

            begin
              gen[59][17].run()  ;
            end
            begin
              drv[59][17].run()  ;
            end
            begin
              dma2mem[59][17].run()  ;
            end

            begin
              gen[59][18].run()  ;
            end
            begin
              drv[59][18].run()  ;
            end
            begin
              dma2mem[59][18].run()  ;
            end

            begin
              gen[59][19].run()  ;
            end
            begin
              drv[59][19].run()  ;
            end
            begin
              dma2mem[59][19].run()  ;
            end

            begin
              gen[59][20].run()  ;
            end
            begin
              drv[59][20].run()  ;
            end
            begin
              dma2mem[59][20].run()  ;
            end

            begin
              gen[59][21].run()  ;
            end
            begin
              drv[59][21].run()  ;
            end
            begin
              dma2mem[59][21].run()  ;
            end

            begin
              gen[59][22].run()  ;
            end
            begin
              drv[59][22].run()  ;
            end
            begin
              dma2mem[59][22].run()  ;
            end

            begin
              gen[59][23].run()  ;
            end
            begin
              drv[59][23].run()  ;
            end
            begin
              dma2mem[59][23].run()  ;
            end

            begin
              gen[59][24].run()  ;
            end
            begin
              drv[59][24].run()  ;
            end
            begin
              dma2mem[59][24].run()  ;
            end

            begin
              gen[59][25].run()  ;
            end
            begin
              drv[59][25].run()  ;
            end
            begin
              dma2mem[59][25].run()  ;
            end

            begin
              gen[59][26].run()  ;
            end
            begin
              drv[59][26].run()  ;
            end
            begin
              dma2mem[59][26].run()  ;
            end

            begin
              gen[59][27].run()  ;
            end
            begin
              drv[59][27].run()  ;
            end
            begin
              dma2mem[59][27].run()  ;
            end

            begin
              gen[59][28].run()  ;
            end
            begin
              drv[59][28].run()  ;
            end
            begin
              dma2mem[59][28].run()  ;
            end

            begin
              gen[59][29].run()  ;
            end
            begin
              drv[59][29].run()  ;
            end
            begin
              dma2mem[59][29].run()  ;
            end

            begin
              gen[59][30].run()  ;
            end
            begin
              drv[59][30].run()  ;
            end
            begin
              dma2mem[59][30].run()  ;
            end

            begin
              gen[59][31].run()  ;
            end
            begin
              drv[59][31].run()  ;
            end
            begin
              dma2mem[59][31].run()  ;
            end

            begin
              gen[60][0].run()  ;
            end
            begin
              drv[60][0].run()  ;
            end
            begin
              dma2mem[60][0].run()  ;
            end

            begin
              gen[60][1].run()  ;
            end
            begin
              drv[60][1].run()  ;
            end
            begin
              dma2mem[60][1].run()  ;
            end

            begin
              gen[60][2].run()  ;
            end
            begin
              drv[60][2].run()  ;
            end
            begin
              dma2mem[60][2].run()  ;
            end

            begin
              gen[60][3].run()  ;
            end
            begin
              drv[60][3].run()  ;
            end
            begin
              dma2mem[60][3].run()  ;
            end

            begin
              gen[60][4].run()  ;
            end
            begin
              drv[60][4].run()  ;
            end
            begin
              dma2mem[60][4].run()  ;
            end

            begin
              gen[60][5].run()  ;
            end
            begin
              drv[60][5].run()  ;
            end
            begin
              dma2mem[60][5].run()  ;
            end

            begin
              gen[60][6].run()  ;
            end
            begin
              drv[60][6].run()  ;
            end
            begin
              dma2mem[60][6].run()  ;
            end

            begin
              gen[60][7].run()  ;
            end
            begin
              drv[60][7].run()  ;
            end
            begin
              dma2mem[60][7].run()  ;
            end

            begin
              gen[60][8].run()  ;
            end
            begin
              drv[60][8].run()  ;
            end
            begin
              dma2mem[60][8].run()  ;
            end

            begin
              gen[60][9].run()  ;
            end
            begin
              drv[60][9].run()  ;
            end
            begin
              dma2mem[60][9].run()  ;
            end

            begin
              gen[60][10].run()  ;
            end
            begin
              drv[60][10].run()  ;
            end
            begin
              dma2mem[60][10].run()  ;
            end

            begin
              gen[60][11].run()  ;
            end
            begin
              drv[60][11].run()  ;
            end
            begin
              dma2mem[60][11].run()  ;
            end

            begin
              gen[60][12].run()  ;
            end
            begin
              drv[60][12].run()  ;
            end
            begin
              dma2mem[60][12].run()  ;
            end

            begin
              gen[60][13].run()  ;
            end
            begin
              drv[60][13].run()  ;
            end
            begin
              dma2mem[60][13].run()  ;
            end

            begin
              gen[60][14].run()  ;
            end
            begin
              drv[60][14].run()  ;
            end
            begin
              dma2mem[60][14].run()  ;
            end

            begin
              gen[60][15].run()  ;
            end
            begin
              drv[60][15].run()  ;
            end
            begin
              dma2mem[60][15].run()  ;
            end

            begin
              gen[60][16].run()  ;
            end
            begin
              drv[60][16].run()  ;
            end
            begin
              dma2mem[60][16].run()  ;
            end

            begin
              gen[60][17].run()  ;
            end
            begin
              drv[60][17].run()  ;
            end
            begin
              dma2mem[60][17].run()  ;
            end

            begin
              gen[60][18].run()  ;
            end
            begin
              drv[60][18].run()  ;
            end
            begin
              dma2mem[60][18].run()  ;
            end

            begin
              gen[60][19].run()  ;
            end
            begin
              drv[60][19].run()  ;
            end
            begin
              dma2mem[60][19].run()  ;
            end

            begin
              gen[60][20].run()  ;
            end
            begin
              drv[60][20].run()  ;
            end
            begin
              dma2mem[60][20].run()  ;
            end

            begin
              gen[60][21].run()  ;
            end
            begin
              drv[60][21].run()  ;
            end
            begin
              dma2mem[60][21].run()  ;
            end

            begin
              gen[60][22].run()  ;
            end
            begin
              drv[60][22].run()  ;
            end
            begin
              dma2mem[60][22].run()  ;
            end

            begin
              gen[60][23].run()  ;
            end
            begin
              drv[60][23].run()  ;
            end
            begin
              dma2mem[60][23].run()  ;
            end

            begin
              gen[60][24].run()  ;
            end
            begin
              drv[60][24].run()  ;
            end
            begin
              dma2mem[60][24].run()  ;
            end

            begin
              gen[60][25].run()  ;
            end
            begin
              drv[60][25].run()  ;
            end
            begin
              dma2mem[60][25].run()  ;
            end

            begin
              gen[60][26].run()  ;
            end
            begin
              drv[60][26].run()  ;
            end
            begin
              dma2mem[60][26].run()  ;
            end

            begin
              gen[60][27].run()  ;
            end
            begin
              drv[60][27].run()  ;
            end
            begin
              dma2mem[60][27].run()  ;
            end

            begin
              gen[60][28].run()  ;
            end
            begin
              drv[60][28].run()  ;
            end
            begin
              dma2mem[60][28].run()  ;
            end

            begin
              gen[60][29].run()  ;
            end
            begin
              drv[60][29].run()  ;
            end
            begin
              dma2mem[60][29].run()  ;
            end

            begin
              gen[60][30].run()  ;
            end
            begin
              drv[60][30].run()  ;
            end
            begin
              dma2mem[60][30].run()  ;
            end

            begin
              gen[60][31].run()  ;
            end
            begin
              drv[60][31].run()  ;
            end
            begin
              dma2mem[60][31].run()  ;
            end

            begin
              gen[61][0].run()  ;
            end
            begin
              drv[61][0].run()  ;
            end
            begin
              dma2mem[61][0].run()  ;
            end

            begin
              gen[61][1].run()  ;
            end
            begin
              drv[61][1].run()  ;
            end
            begin
              dma2mem[61][1].run()  ;
            end

            begin
              gen[61][2].run()  ;
            end
            begin
              drv[61][2].run()  ;
            end
            begin
              dma2mem[61][2].run()  ;
            end

            begin
              gen[61][3].run()  ;
            end
            begin
              drv[61][3].run()  ;
            end
            begin
              dma2mem[61][3].run()  ;
            end

            begin
              gen[61][4].run()  ;
            end
            begin
              drv[61][4].run()  ;
            end
            begin
              dma2mem[61][4].run()  ;
            end

            begin
              gen[61][5].run()  ;
            end
            begin
              drv[61][5].run()  ;
            end
            begin
              dma2mem[61][5].run()  ;
            end

            begin
              gen[61][6].run()  ;
            end
            begin
              drv[61][6].run()  ;
            end
            begin
              dma2mem[61][6].run()  ;
            end

            begin
              gen[61][7].run()  ;
            end
            begin
              drv[61][7].run()  ;
            end
            begin
              dma2mem[61][7].run()  ;
            end

            begin
              gen[61][8].run()  ;
            end
            begin
              drv[61][8].run()  ;
            end
            begin
              dma2mem[61][8].run()  ;
            end

            begin
              gen[61][9].run()  ;
            end
            begin
              drv[61][9].run()  ;
            end
            begin
              dma2mem[61][9].run()  ;
            end

            begin
              gen[61][10].run()  ;
            end
            begin
              drv[61][10].run()  ;
            end
            begin
              dma2mem[61][10].run()  ;
            end

            begin
              gen[61][11].run()  ;
            end
            begin
              drv[61][11].run()  ;
            end
            begin
              dma2mem[61][11].run()  ;
            end

            begin
              gen[61][12].run()  ;
            end
            begin
              drv[61][12].run()  ;
            end
            begin
              dma2mem[61][12].run()  ;
            end

            begin
              gen[61][13].run()  ;
            end
            begin
              drv[61][13].run()  ;
            end
            begin
              dma2mem[61][13].run()  ;
            end

            begin
              gen[61][14].run()  ;
            end
            begin
              drv[61][14].run()  ;
            end
            begin
              dma2mem[61][14].run()  ;
            end

            begin
              gen[61][15].run()  ;
            end
            begin
              drv[61][15].run()  ;
            end
            begin
              dma2mem[61][15].run()  ;
            end

            begin
              gen[61][16].run()  ;
            end
            begin
              drv[61][16].run()  ;
            end
            begin
              dma2mem[61][16].run()  ;
            end

            begin
              gen[61][17].run()  ;
            end
            begin
              drv[61][17].run()  ;
            end
            begin
              dma2mem[61][17].run()  ;
            end

            begin
              gen[61][18].run()  ;
            end
            begin
              drv[61][18].run()  ;
            end
            begin
              dma2mem[61][18].run()  ;
            end

            begin
              gen[61][19].run()  ;
            end
            begin
              drv[61][19].run()  ;
            end
            begin
              dma2mem[61][19].run()  ;
            end

            begin
              gen[61][20].run()  ;
            end
            begin
              drv[61][20].run()  ;
            end
            begin
              dma2mem[61][20].run()  ;
            end

            begin
              gen[61][21].run()  ;
            end
            begin
              drv[61][21].run()  ;
            end
            begin
              dma2mem[61][21].run()  ;
            end

            begin
              gen[61][22].run()  ;
            end
            begin
              drv[61][22].run()  ;
            end
            begin
              dma2mem[61][22].run()  ;
            end

            begin
              gen[61][23].run()  ;
            end
            begin
              drv[61][23].run()  ;
            end
            begin
              dma2mem[61][23].run()  ;
            end

            begin
              gen[61][24].run()  ;
            end
            begin
              drv[61][24].run()  ;
            end
            begin
              dma2mem[61][24].run()  ;
            end

            begin
              gen[61][25].run()  ;
            end
            begin
              drv[61][25].run()  ;
            end
            begin
              dma2mem[61][25].run()  ;
            end

            begin
              gen[61][26].run()  ;
            end
            begin
              drv[61][26].run()  ;
            end
            begin
              dma2mem[61][26].run()  ;
            end

            begin
              gen[61][27].run()  ;
            end
            begin
              drv[61][27].run()  ;
            end
            begin
              dma2mem[61][27].run()  ;
            end

            begin
              gen[61][28].run()  ;
            end
            begin
              drv[61][28].run()  ;
            end
            begin
              dma2mem[61][28].run()  ;
            end

            begin
              gen[61][29].run()  ;
            end
            begin
              drv[61][29].run()  ;
            end
            begin
              dma2mem[61][29].run()  ;
            end

            begin
              gen[61][30].run()  ;
            end
            begin
              drv[61][30].run()  ;
            end
            begin
              dma2mem[61][30].run()  ;
            end

            begin
              gen[61][31].run()  ;
            end
            begin
              drv[61][31].run()  ;
            end
            begin
              dma2mem[61][31].run()  ;
            end

            begin
              gen[62][0].run()  ;
            end
            begin
              drv[62][0].run()  ;
            end
            begin
              dma2mem[62][0].run()  ;
            end

            begin
              gen[62][1].run()  ;
            end
            begin
              drv[62][1].run()  ;
            end
            begin
              dma2mem[62][1].run()  ;
            end

            begin
              gen[62][2].run()  ;
            end
            begin
              drv[62][2].run()  ;
            end
            begin
              dma2mem[62][2].run()  ;
            end

            begin
              gen[62][3].run()  ;
            end
            begin
              drv[62][3].run()  ;
            end
            begin
              dma2mem[62][3].run()  ;
            end

            begin
              gen[62][4].run()  ;
            end
            begin
              drv[62][4].run()  ;
            end
            begin
              dma2mem[62][4].run()  ;
            end

            begin
              gen[62][5].run()  ;
            end
            begin
              drv[62][5].run()  ;
            end
            begin
              dma2mem[62][5].run()  ;
            end

            begin
              gen[62][6].run()  ;
            end
            begin
              drv[62][6].run()  ;
            end
            begin
              dma2mem[62][6].run()  ;
            end

            begin
              gen[62][7].run()  ;
            end
            begin
              drv[62][7].run()  ;
            end
            begin
              dma2mem[62][7].run()  ;
            end

            begin
              gen[62][8].run()  ;
            end
            begin
              drv[62][8].run()  ;
            end
            begin
              dma2mem[62][8].run()  ;
            end

            begin
              gen[62][9].run()  ;
            end
            begin
              drv[62][9].run()  ;
            end
            begin
              dma2mem[62][9].run()  ;
            end

            begin
              gen[62][10].run()  ;
            end
            begin
              drv[62][10].run()  ;
            end
            begin
              dma2mem[62][10].run()  ;
            end

            begin
              gen[62][11].run()  ;
            end
            begin
              drv[62][11].run()  ;
            end
            begin
              dma2mem[62][11].run()  ;
            end

            begin
              gen[62][12].run()  ;
            end
            begin
              drv[62][12].run()  ;
            end
            begin
              dma2mem[62][12].run()  ;
            end

            begin
              gen[62][13].run()  ;
            end
            begin
              drv[62][13].run()  ;
            end
            begin
              dma2mem[62][13].run()  ;
            end

            begin
              gen[62][14].run()  ;
            end
            begin
              drv[62][14].run()  ;
            end
            begin
              dma2mem[62][14].run()  ;
            end

            begin
              gen[62][15].run()  ;
            end
            begin
              drv[62][15].run()  ;
            end
            begin
              dma2mem[62][15].run()  ;
            end

            begin
              gen[62][16].run()  ;
            end
            begin
              drv[62][16].run()  ;
            end
            begin
              dma2mem[62][16].run()  ;
            end

            begin
              gen[62][17].run()  ;
            end
            begin
              drv[62][17].run()  ;
            end
            begin
              dma2mem[62][17].run()  ;
            end

            begin
              gen[62][18].run()  ;
            end
            begin
              drv[62][18].run()  ;
            end
            begin
              dma2mem[62][18].run()  ;
            end

            begin
              gen[62][19].run()  ;
            end
            begin
              drv[62][19].run()  ;
            end
            begin
              dma2mem[62][19].run()  ;
            end

            begin
              gen[62][20].run()  ;
            end
            begin
              drv[62][20].run()  ;
            end
            begin
              dma2mem[62][20].run()  ;
            end

            begin
              gen[62][21].run()  ;
            end
            begin
              drv[62][21].run()  ;
            end
            begin
              dma2mem[62][21].run()  ;
            end

            begin
              gen[62][22].run()  ;
            end
            begin
              drv[62][22].run()  ;
            end
            begin
              dma2mem[62][22].run()  ;
            end

            begin
              gen[62][23].run()  ;
            end
            begin
              drv[62][23].run()  ;
            end
            begin
              dma2mem[62][23].run()  ;
            end

            begin
              gen[62][24].run()  ;
            end
            begin
              drv[62][24].run()  ;
            end
            begin
              dma2mem[62][24].run()  ;
            end

            begin
              gen[62][25].run()  ;
            end
            begin
              drv[62][25].run()  ;
            end
            begin
              dma2mem[62][25].run()  ;
            end

            begin
              gen[62][26].run()  ;
            end
            begin
              drv[62][26].run()  ;
            end
            begin
              dma2mem[62][26].run()  ;
            end

            begin
              gen[62][27].run()  ;
            end
            begin
              drv[62][27].run()  ;
            end
            begin
              dma2mem[62][27].run()  ;
            end

            begin
              gen[62][28].run()  ;
            end
            begin
              drv[62][28].run()  ;
            end
            begin
              dma2mem[62][28].run()  ;
            end

            begin
              gen[62][29].run()  ;
            end
            begin
              drv[62][29].run()  ;
            end
            begin
              dma2mem[62][29].run()  ;
            end

            begin
              gen[62][30].run()  ;
            end
            begin
              drv[62][30].run()  ;
            end
            begin
              dma2mem[62][30].run()  ;
            end

            begin
              gen[62][31].run()  ;
            end
            begin
              drv[62][31].run()  ;
            end
            begin
              dma2mem[62][31].run()  ;
            end

            begin
              gen[63][0].run()  ;
            end
            begin
              drv[63][0].run()  ;
            end
            begin
              dma2mem[63][0].run()  ;
            end

            begin
              gen[63][1].run()  ;
            end
            begin
              drv[63][1].run()  ;
            end
            begin
              dma2mem[63][1].run()  ;
            end

            begin
              gen[63][2].run()  ;
            end
            begin
              drv[63][2].run()  ;
            end
            begin
              dma2mem[63][2].run()  ;
            end

            begin
              gen[63][3].run()  ;
            end
            begin
              drv[63][3].run()  ;
            end
            begin
              dma2mem[63][3].run()  ;
            end

            begin
              gen[63][4].run()  ;
            end
            begin
              drv[63][4].run()  ;
            end
            begin
              dma2mem[63][4].run()  ;
            end

            begin
              gen[63][5].run()  ;
            end
            begin
              drv[63][5].run()  ;
            end
            begin
              dma2mem[63][5].run()  ;
            end

            begin
              gen[63][6].run()  ;
            end
            begin
              drv[63][6].run()  ;
            end
            begin
              dma2mem[63][6].run()  ;
            end

            begin
              gen[63][7].run()  ;
            end
            begin
              drv[63][7].run()  ;
            end
            begin
              dma2mem[63][7].run()  ;
            end

            begin
              gen[63][8].run()  ;
            end
            begin
              drv[63][8].run()  ;
            end
            begin
              dma2mem[63][8].run()  ;
            end

            begin
              gen[63][9].run()  ;
            end
            begin
              drv[63][9].run()  ;
            end
            begin
              dma2mem[63][9].run()  ;
            end

            begin
              gen[63][10].run()  ;
            end
            begin
              drv[63][10].run()  ;
            end
            begin
              dma2mem[63][10].run()  ;
            end

            begin
              gen[63][11].run()  ;
            end
            begin
              drv[63][11].run()  ;
            end
            begin
              dma2mem[63][11].run()  ;
            end

            begin
              gen[63][12].run()  ;
            end
            begin
              drv[63][12].run()  ;
            end
            begin
              dma2mem[63][12].run()  ;
            end

            begin
              gen[63][13].run()  ;
            end
            begin
              drv[63][13].run()  ;
            end
            begin
              dma2mem[63][13].run()  ;
            end

            begin
              gen[63][14].run()  ;
            end
            begin
              drv[63][14].run()  ;
            end
            begin
              dma2mem[63][14].run()  ;
            end

            begin
              gen[63][15].run()  ;
            end
            begin
              drv[63][15].run()  ;
            end
            begin
              dma2mem[63][15].run()  ;
            end

            begin
              gen[63][16].run()  ;
            end
            begin
              drv[63][16].run()  ;
            end
            begin
              dma2mem[63][16].run()  ;
            end

            begin
              gen[63][17].run()  ;
            end
            begin
              drv[63][17].run()  ;
            end
            begin
              dma2mem[63][17].run()  ;
            end

            begin
              gen[63][18].run()  ;
            end
            begin
              drv[63][18].run()  ;
            end
            begin
              dma2mem[63][18].run()  ;
            end

            begin
              gen[63][19].run()  ;
            end
            begin
              drv[63][19].run()  ;
            end
            begin
              dma2mem[63][19].run()  ;
            end

            begin
              gen[63][20].run()  ;
            end
            begin
              drv[63][20].run()  ;
            end
            begin
              dma2mem[63][20].run()  ;
            end

            begin
              gen[63][21].run()  ;
            end
            begin
              drv[63][21].run()  ;
            end
            begin
              dma2mem[63][21].run()  ;
            end

            begin
              gen[63][22].run()  ;
            end
            begin
              drv[63][22].run()  ;
            end
            begin
              dma2mem[63][22].run()  ;
            end

            begin
              gen[63][23].run()  ;
            end
            begin
              drv[63][23].run()  ;
            end
            begin
              dma2mem[63][23].run()  ;
            end

            begin
              gen[63][24].run()  ;
            end
            begin
              drv[63][24].run()  ;
            end
            begin
              dma2mem[63][24].run()  ;
            end

            begin
              gen[63][25].run()  ;
            end
            begin
              drv[63][25].run()  ;
            end
            begin
              dma2mem[63][25].run()  ;
            end

            begin
              gen[63][26].run()  ;
            end
            begin
              drv[63][26].run()  ;
            end
            begin
              dma2mem[63][26].run()  ;
            end

            begin
              gen[63][27].run()  ;
            end
            begin
              drv[63][27].run()  ;
            end
            begin
              dma2mem[63][27].run()  ;
            end

            begin
              gen[63][28].run()  ;
            end
            begin
              drv[63][28].run()  ;
            end
            begin
              dma2mem[63][28].run()  ;
            end

            begin
              gen[63][29].run()  ;
            end
            begin
              drv[63][29].run()  ;
            end
            begin
              dma2mem[63][29].run()  ;
            end

            begin
              gen[63][30].run()  ;
            end
            begin
              drv[63][30].run()  ;
            end
            begin
              dma2mem[63][30].run()  ;
            end

            begin
              gen[63][31].run()  ;
            end
            begin
              drv[63][31].run()  ;
            end
            begin
              dma2mem[63][31].run()  ;
            end
