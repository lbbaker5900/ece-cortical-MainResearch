
  // Lane 0, Stream 0
  wire                                         sdp__std__lane0_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane0_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane0_strm0_data          ;
  wire                                         std__sdp__lane0_strm0_data_valid    ;
  // Lane 1, Stream 0
  wire                                         sdp__std__lane1_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane1_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane1_strm0_data          ;
  wire                                         std__sdp__lane1_strm0_data_valid    ;
  // Lane 2, Stream 0
  wire                                         sdp__std__lane2_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane2_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane2_strm0_data          ;
  wire                                         std__sdp__lane2_strm0_data_valid    ;
  // Lane 3, Stream 0
  wire                                         sdp__std__lane3_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane3_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane3_strm0_data          ;
  wire                                         std__sdp__lane3_strm0_data_valid    ;
  // Lane 4, Stream 0
  wire                                         sdp__std__lane4_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane4_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane4_strm0_data          ;
  wire                                         std__sdp__lane4_strm0_data_valid    ;
  // Lane 5, Stream 0
  wire                                         sdp__std__lane5_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane5_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane5_strm0_data          ;
  wire                                         std__sdp__lane5_strm0_data_valid    ;
  // Lane 6, Stream 0
  wire                                         sdp__std__lane6_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane6_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane6_strm0_data          ;
  wire                                         std__sdp__lane6_strm0_data_valid    ;
  // Lane 7, Stream 0
  wire                                         sdp__std__lane7_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane7_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane7_strm0_data          ;
  wire                                         std__sdp__lane7_strm0_data_valid    ;
  // Lane 8, Stream 0
  wire                                         sdp__std__lane8_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane8_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane8_strm0_data          ;
  wire                                         std__sdp__lane8_strm0_data_valid    ;
  // Lane 9, Stream 0
  wire                                         sdp__std__lane9_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane9_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane9_strm0_data          ;
  wire                                         std__sdp__lane9_strm0_data_valid    ;
  // Lane 10, Stream 0
  wire                                         sdp__std__lane10_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane10_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane10_strm0_data          ;
  wire                                         std__sdp__lane10_strm0_data_valid    ;
  // Lane 11, Stream 0
  wire                                         sdp__std__lane11_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane11_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane11_strm0_data          ;
  wire                                         std__sdp__lane11_strm0_data_valid    ;
  // Lane 12, Stream 0
  wire                                         sdp__std__lane12_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane12_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane12_strm0_data          ;
  wire                                         std__sdp__lane12_strm0_data_valid    ;
  // Lane 13, Stream 0
  wire                                         sdp__std__lane13_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane13_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane13_strm0_data          ;
  wire                                         std__sdp__lane13_strm0_data_valid    ;
  // Lane 14, Stream 0
  wire                                         sdp__std__lane14_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane14_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane14_strm0_data          ;
  wire                                         std__sdp__lane14_strm0_data_valid    ;
  // Lane 15, Stream 0
  wire                                         sdp__std__lane15_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane15_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane15_strm0_data          ;
  wire                                         std__sdp__lane15_strm0_data_valid    ;
  // Lane 16, Stream 0
  wire                                         sdp__std__lane16_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane16_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane16_strm0_data          ;
  wire                                         std__sdp__lane16_strm0_data_valid    ;
  // Lane 17, Stream 0
  wire                                         sdp__std__lane17_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane17_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane17_strm0_data          ;
  wire                                         std__sdp__lane17_strm0_data_valid    ;
  // Lane 18, Stream 0
  wire                                         sdp__std__lane18_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane18_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane18_strm0_data          ;
  wire                                         std__sdp__lane18_strm0_data_valid    ;
  // Lane 19, Stream 0
  wire                                         sdp__std__lane19_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane19_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane19_strm0_data          ;
  wire                                         std__sdp__lane19_strm0_data_valid    ;
  // Lane 20, Stream 0
  wire                                         sdp__std__lane20_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane20_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane20_strm0_data          ;
  wire                                         std__sdp__lane20_strm0_data_valid    ;
  // Lane 21, Stream 0
  wire                                         sdp__std__lane21_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane21_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane21_strm0_data          ;
  wire                                         std__sdp__lane21_strm0_data_valid    ;
  // Lane 22, Stream 0
  wire                                         sdp__std__lane22_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane22_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane22_strm0_data          ;
  wire                                         std__sdp__lane22_strm0_data_valid    ;
  // Lane 23, Stream 0
  wire                                         sdp__std__lane23_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane23_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane23_strm0_data          ;
  wire                                         std__sdp__lane23_strm0_data_valid    ;
  // Lane 24, Stream 0
  wire                                         sdp__std__lane24_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane24_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane24_strm0_data          ;
  wire                                         std__sdp__lane24_strm0_data_valid    ;
  // Lane 25, Stream 0
  wire                                         sdp__std__lane25_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane25_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane25_strm0_data          ;
  wire                                         std__sdp__lane25_strm0_data_valid    ;
  // Lane 26, Stream 0
  wire                                         sdp__std__lane26_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane26_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane26_strm0_data          ;
  wire                                         std__sdp__lane26_strm0_data_valid    ;
  // Lane 27, Stream 0
  wire                                         sdp__std__lane27_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane27_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane27_strm0_data          ;
  wire                                         std__sdp__lane27_strm0_data_valid    ;
  // Lane 28, Stream 0
  wire                                         sdp__std__lane28_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane28_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane28_strm0_data          ;
  wire                                         std__sdp__lane28_strm0_data_valid    ;
  // Lane 29, Stream 0
  wire                                         sdp__std__lane29_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane29_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane29_strm0_data          ;
  wire                                         std__sdp__lane29_strm0_data_valid    ;
  // Lane 30, Stream 0
  wire                                         sdp__std__lane30_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane30_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane30_strm0_data          ;
  wire                                         std__sdp__lane30_strm0_data_valid    ;
  // Lane 31, Stream 0
  wire                                         sdp__std__lane31_strm0_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane31_strm0_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane31_strm0_data          ;
  wire                                         std__sdp__lane31_strm0_data_valid    ;

  // Lane 0, Stream 1
  wire                                         sdp__std__lane0_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane0_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane0_strm1_data          ;
  wire                                         std__sdp__lane0_strm1_data_valid    ;
  // Lane 1, Stream 1
  wire                                         sdp__std__lane1_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane1_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane1_strm1_data          ;
  wire                                         std__sdp__lane1_strm1_data_valid    ;
  // Lane 2, Stream 1
  wire                                         sdp__std__lane2_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane2_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane2_strm1_data          ;
  wire                                         std__sdp__lane2_strm1_data_valid    ;
  // Lane 3, Stream 1
  wire                                         sdp__std__lane3_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane3_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane3_strm1_data          ;
  wire                                         std__sdp__lane3_strm1_data_valid    ;
  // Lane 4, Stream 1
  wire                                         sdp__std__lane4_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane4_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane4_strm1_data          ;
  wire                                         std__sdp__lane4_strm1_data_valid    ;
  // Lane 5, Stream 1
  wire                                         sdp__std__lane5_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane5_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane5_strm1_data          ;
  wire                                         std__sdp__lane5_strm1_data_valid    ;
  // Lane 6, Stream 1
  wire                                         sdp__std__lane6_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane6_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane6_strm1_data          ;
  wire                                         std__sdp__lane6_strm1_data_valid    ;
  // Lane 7, Stream 1
  wire                                         sdp__std__lane7_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane7_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane7_strm1_data          ;
  wire                                         std__sdp__lane7_strm1_data_valid    ;
  // Lane 8, Stream 1
  wire                                         sdp__std__lane8_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane8_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane8_strm1_data          ;
  wire                                         std__sdp__lane8_strm1_data_valid    ;
  // Lane 9, Stream 1
  wire                                         sdp__std__lane9_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane9_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane9_strm1_data          ;
  wire                                         std__sdp__lane9_strm1_data_valid    ;
  // Lane 10, Stream 1
  wire                                         sdp__std__lane10_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane10_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane10_strm1_data          ;
  wire                                         std__sdp__lane10_strm1_data_valid    ;
  // Lane 11, Stream 1
  wire                                         sdp__std__lane11_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane11_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane11_strm1_data          ;
  wire                                         std__sdp__lane11_strm1_data_valid    ;
  // Lane 12, Stream 1
  wire                                         sdp__std__lane12_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane12_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane12_strm1_data          ;
  wire                                         std__sdp__lane12_strm1_data_valid    ;
  // Lane 13, Stream 1
  wire                                         sdp__std__lane13_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane13_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane13_strm1_data          ;
  wire                                         std__sdp__lane13_strm1_data_valid    ;
  // Lane 14, Stream 1
  wire                                         sdp__std__lane14_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane14_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane14_strm1_data          ;
  wire                                         std__sdp__lane14_strm1_data_valid    ;
  // Lane 15, Stream 1
  wire                                         sdp__std__lane15_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane15_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane15_strm1_data          ;
  wire                                         std__sdp__lane15_strm1_data_valid    ;
  // Lane 16, Stream 1
  wire                                         sdp__std__lane16_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane16_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane16_strm1_data          ;
  wire                                         std__sdp__lane16_strm1_data_valid    ;
  // Lane 17, Stream 1
  wire                                         sdp__std__lane17_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane17_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane17_strm1_data          ;
  wire                                         std__sdp__lane17_strm1_data_valid    ;
  // Lane 18, Stream 1
  wire                                         sdp__std__lane18_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane18_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane18_strm1_data          ;
  wire                                         std__sdp__lane18_strm1_data_valid    ;
  // Lane 19, Stream 1
  wire                                         sdp__std__lane19_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane19_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane19_strm1_data          ;
  wire                                         std__sdp__lane19_strm1_data_valid    ;
  // Lane 20, Stream 1
  wire                                         sdp__std__lane20_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane20_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane20_strm1_data          ;
  wire                                         std__sdp__lane20_strm1_data_valid    ;
  // Lane 21, Stream 1
  wire                                         sdp__std__lane21_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane21_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane21_strm1_data          ;
  wire                                         std__sdp__lane21_strm1_data_valid    ;
  // Lane 22, Stream 1
  wire                                         sdp__std__lane22_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane22_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane22_strm1_data          ;
  wire                                         std__sdp__lane22_strm1_data_valid    ;
  // Lane 23, Stream 1
  wire                                         sdp__std__lane23_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane23_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane23_strm1_data          ;
  wire                                         std__sdp__lane23_strm1_data_valid    ;
  // Lane 24, Stream 1
  wire                                         sdp__std__lane24_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane24_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane24_strm1_data          ;
  wire                                         std__sdp__lane24_strm1_data_valid    ;
  // Lane 25, Stream 1
  wire                                         sdp__std__lane25_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane25_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane25_strm1_data          ;
  wire                                         std__sdp__lane25_strm1_data_valid    ;
  // Lane 26, Stream 1
  wire                                         sdp__std__lane26_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane26_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane26_strm1_data          ;
  wire                                         std__sdp__lane26_strm1_data_valid    ;
  // Lane 27, Stream 1
  wire                                         sdp__std__lane27_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane27_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane27_strm1_data          ;
  wire                                         std__sdp__lane27_strm1_data_valid    ;
  // Lane 28, Stream 1
  wire                                         sdp__std__lane28_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane28_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane28_strm1_data          ;
  wire                                         std__sdp__lane28_strm1_data_valid    ;
  // Lane 29, Stream 1
  wire                                         sdp__std__lane29_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane29_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane29_strm1_data          ;
  wire                                         std__sdp__lane29_strm1_data_valid    ;
  // Lane 30, Stream 1
  wire                                         sdp__std__lane30_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane30_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane30_strm1_data          ;
  wire                                         std__sdp__lane30_strm1_data_valid    ;
  // Lane 31, Stream 1
  wire                                         sdp__std__lane31_strm1_ready         ;
  wire  [`DMA_CONT_STRM_CNTL_RANGE     ]       std__sdp__lane31_strm1_cntl          ;
  wire  [`STREAMING_OP_DATA_RANGE      ]       std__sdp__lane31_strm1_data          ;
  wire                                         std__sdp__lane31_strm1_data_valid    ;
