
  input                                             stOp__sti__lane0_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane0_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane0_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane0_strm0_data_mask   ;
  output                                            sti__stOp__lane0_strm0_data_valid  ;

  input                                             stOp__sti__lane0_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane0_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane0_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane0_strm1_data_mask   ;
  output                                            sti__stOp__lane0_strm1_data_valid  ;

  input                                             stOp__sti__lane1_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane1_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane1_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane1_strm0_data_mask   ;
  output                                            sti__stOp__lane1_strm0_data_valid  ;

  input                                             stOp__sti__lane1_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane1_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane1_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane1_strm1_data_mask   ;
  output                                            sti__stOp__lane1_strm1_data_valid  ;

  input                                             stOp__sti__lane2_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane2_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane2_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane2_strm0_data_mask   ;
  output                                            sti__stOp__lane2_strm0_data_valid  ;

  input                                             stOp__sti__lane2_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane2_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane2_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane2_strm1_data_mask   ;
  output                                            sti__stOp__lane2_strm1_data_valid  ;

  input                                             stOp__sti__lane3_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane3_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane3_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane3_strm0_data_mask   ;
  output                                            sti__stOp__lane3_strm0_data_valid  ;

  input                                             stOp__sti__lane3_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane3_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane3_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane3_strm1_data_mask   ;
  output                                            sti__stOp__lane3_strm1_data_valid  ;

  input                                             stOp__sti__lane4_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane4_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane4_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane4_strm0_data_mask   ;
  output                                            sti__stOp__lane4_strm0_data_valid  ;

  input                                             stOp__sti__lane4_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane4_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane4_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane4_strm1_data_mask   ;
  output                                            sti__stOp__lane4_strm1_data_valid  ;

  input                                             stOp__sti__lane5_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane5_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane5_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane5_strm0_data_mask   ;
  output                                            sti__stOp__lane5_strm0_data_valid  ;

  input                                             stOp__sti__lane5_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane5_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane5_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane5_strm1_data_mask   ;
  output                                            sti__stOp__lane5_strm1_data_valid  ;

  input                                             stOp__sti__lane6_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane6_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane6_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane6_strm0_data_mask   ;
  output                                            sti__stOp__lane6_strm0_data_valid  ;

  input                                             stOp__sti__lane6_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane6_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane6_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane6_strm1_data_mask   ;
  output                                            sti__stOp__lane6_strm1_data_valid  ;

  input                                             stOp__sti__lane7_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane7_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane7_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane7_strm0_data_mask   ;
  output                                            sti__stOp__lane7_strm0_data_valid  ;

  input                                             stOp__sti__lane7_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane7_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane7_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane7_strm1_data_mask   ;
  output                                            sti__stOp__lane7_strm1_data_valid  ;

  input                                             stOp__sti__lane8_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane8_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane8_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane8_strm0_data_mask   ;
  output                                            sti__stOp__lane8_strm0_data_valid  ;

  input                                             stOp__sti__lane8_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane8_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane8_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane8_strm1_data_mask   ;
  output                                            sti__stOp__lane8_strm1_data_valid  ;

  input                                             stOp__sti__lane9_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane9_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane9_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane9_strm0_data_mask   ;
  output                                            sti__stOp__lane9_strm0_data_valid  ;

  input                                             stOp__sti__lane9_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane9_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane9_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane9_strm1_data_mask   ;
  output                                            sti__stOp__lane9_strm1_data_valid  ;

  input                                             stOp__sti__lane10_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane10_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane10_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane10_strm0_data_mask   ;
  output                                            sti__stOp__lane10_strm0_data_valid  ;

  input                                             stOp__sti__lane10_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane10_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane10_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane10_strm1_data_mask   ;
  output                                            sti__stOp__lane10_strm1_data_valid  ;

  input                                             stOp__sti__lane11_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane11_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane11_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane11_strm0_data_mask   ;
  output                                            sti__stOp__lane11_strm0_data_valid  ;

  input                                             stOp__sti__lane11_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane11_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane11_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane11_strm1_data_mask   ;
  output                                            sti__stOp__lane11_strm1_data_valid  ;

  input                                             stOp__sti__lane12_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane12_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane12_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane12_strm0_data_mask   ;
  output                                            sti__stOp__lane12_strm0_data_valid  ;

  input                                             stOp__sti__lane12_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane12_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane12_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane12_strm1_data_mask   ;
  output                                            sti__stOp__lane12_strm1_data_valid  ;

  input                                             stOp__sti__lane13_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane13_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane13_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane13_strm0_data_mask   ;
  output                                            sti__stOp__lane13_strm0_data_valid  ;

  input                                             stOp__sti__lane13_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane13_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane13_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane13_strm1_data_mask   ;
  output                                            sti__stOp__lane13_strm1_data_valid  ;

  input                                             stOp__sti__lane14_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane14_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane14_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane14_strm0_data_mask   ;
  output                                            sti__stOp__lane14_strm0_data_valid  ;

  input                                             stOp__sti__lane14_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane14_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane14_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane14_strm1_data_mask   ;
  output                                            sti__stOp__lane14_strm1_data_valid  ;

  input                                             stOp__sti__lane15_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane15_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane15_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane15_strm0_data_mask   ;
  output                                            sti__stOp__lane15_strm0_data_valid  ;

  input                                             stOp__sti__lane15_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane15_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane15_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane15_strm1_data_mask   ;
  output                                            sti__stOp__lane15_strm1_data_valid  ;

  input                                             stOp__sti__lane16_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane16_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane16_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane16_strm0_data_mask   ;
  output                                            sti__stOp__lane16_strm0_data_valid  ;

  input                                             stOp__sti__lane16_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane16_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane16_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane16_strm1_data_mask   ;
  output                                            sti__stOp__lane16_strm1_data_valid  ;

  input                                             stOp__sti__lane17_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane17_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane17_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane17_strm0_data_mask   ;
  output                                            sti__stOp__lane17_strm0_data_valid  ;

  input                                             stOp__sti__lane17_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane17_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane17_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane17_strm1_data_mask   ;
  output                                            sti__stOp__lane17_strm1_data_valid  ;

  input                                             stOp__sti__lane18_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane18_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane18_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane18_strm0_data_mask   ;
  output                                            sti__stOp__lane18_strm0_data_valid  ;

  input                                             stOp__sti__lane18_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane18_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane18_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane18_strm1_data_mask   ;
  output                                            sti__stOp__lane18_strm1_data_valid  ;

  input                                             stOp__sti__lane19_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane19_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane19_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane19_strm0_data_mask   ;
  output                                            sti__stOp__lane19_strm0_data_valid  ;

  input                                             stOp__sti__lane19_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane19_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane19_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane19_strm1_data_mask   ;
  output                                            sti__stOp__lane19_strm1_data_valid  ;

  input                                             stOp__sti__lane20_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane20_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane20_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane20_strm0_data_mask   ;
  output                                            sti__stOp__lane20_strm0_data_valid  ;

  input                                             stOp__sti__lane20_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane20_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane20_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane20_strm1_data_mask   ;
  output                                            sti__stOp__lane20_strm1_data_valid  ;

  input                                             stOp__sti__lane21_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane21_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane21_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane21_strm0_data_mask   ;
  output                                            sti__stOp__lane21_strm0_data_valid  ;

  input                                             stOp__sti__lane21_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane21_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane21_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane21_strm1_data_mask   ;
  output                                            sti__stOp__lane21_strm1_data_valid  ;

  input                                             stOp__sti__lane22_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane22_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane22_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane22_strm0_data_mask   ;
  output                                            sti__stOp__lane22_strm0_data_valid  ;

  input                                             stOp__sti__lane22_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane22_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane22_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane22_strm1_data_mask   ;
  output                                            sti__stOp__lane22_strm1_data_valid  ;

  input                                             stOp__sti__lane23_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane23_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane23_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane23_strm0_data_mask   ;
  output                                            sti__stOp__lane23_strm0_data_valid  ;

  input                                             stOp__sti__lane23_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane23_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane23_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane23_strm1_data_mask   ;
  output                                            sti__stOp__lane23_strm1_data_valid  ;

  input                                             stOp__sti__lane24_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane24_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane24_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane24_strm0_data_mask   ;
  output                                            sti__stOp__lane24_strm0_data_valid  ;

  input                                             stOp__sti__lane24_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane24_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane24_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane24_strm1_data_mask   ;
  output                                            sti__stOp__lane24_strm1_data_valid  ;

  input                                             stOp__sti__lane25_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane25_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane25_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane25_strm0_data_mask   ;
  output                                            sti__stOp__lane25_strm0_data_valid  ;

  input                                             stOp__sti__lane25_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane25_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane25_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane25_strm1_data_mask   ;
  output                                            sti__stOp__lane25_strm1_data_valid  ;

  input                                             stOp__sti__lane26_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane26_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane26_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane26_strm0_data_mask   ;
  output                                            sti__stOp__lane26_strm0_data_valid  ;

  input                                             stOp__sti__lane26_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane26_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane26_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane26_strm1_data_mask   ;
  output                                            sti__stOp__lane26_strm1_data_valid  ;

  input                                             stOp__sti__lane27_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane27_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane27_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane27_strm0_data_mask   ;
  output                                            sti__stOp__lane27_strm0_data_valid  ;

  input                                             stOp__sti__lane27_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane27_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane27_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane27_strm1_data_mask   ;
  output                                            sti__stOp__lane27_strm1_data_valid  ;

  input                                             stOp__sti__lane28_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane28_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane28_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane28_strm0_data_mask   ;
  output                                            sti__stOp__lane28_strm0_data_valid  ;

  input                                             stOp__sti__lane28_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane28_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane28_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane28_strm1_data_mask   ;
  output                                            sti__stOp__lane28_strm1_data_valid  ;

  input                                             stOp__sti__lane29_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane29_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane29_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane29_strm0_data_mask   ;
  output                                            sti__stOp__lane29_strm0_data_valid  ;

  input                                             stOp__sti__lane29_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane29_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane29_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane29_strm1_data_mask   ;
  output                                            sti__stOp__lane29_strm1_data_valid  ;

  input                                             stOp__sti__lane30_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane30_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane30_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane30_strm0_data_mask   ;
  output                                            sti__stOp__lane30_strm0_data_valid  ;

  input                                             stOp__sti__lane30_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane30_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane30_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane30_strm1_data_mask   ;
  output                                            sti__stOp__lane30_strm1_data_valid  ;

  input                                             stOp__sti__lane31_strm0_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane31_strm0_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane31_strm0_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane31_strm0_data_mask   ;
  output                                            sti__stOp__lane31_strm0_data_valid  ;

  input                                             stOp__sti__lane31_strm1_ready       ;
  output [`COMMON_STD_INTF_CNTL_RANGE       ]       sti__stOp__lane31_strm1_cntl        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane31_strm1_data        ;
  output [`STACK_DOWN_INTF_STRM_DATA_RANGE  ]       sti__stOp__lane31_strm1_data_mask   ;
  output                                            sti__stOp__lane31_strm1_data_valid  ;
