
                  //----------------------------------------------------------------------------------------------------
                  // PE 0
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[0][0].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[0][0].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[0][0].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[0][0].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[0][0].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[0][0].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[0][0].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[0][0].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[0][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[0][0].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[0][1].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[0][1].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[0][1].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[0][1].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[0][1].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[0][1].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[0][1].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[0][1].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[0][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[0][1].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[0][2].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[0][2].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[0][2].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[0][2].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[0][2].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[0][2].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[0][2].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[0][2].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[0][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[0][2].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[0][3].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[0][3].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[0][3].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[0][3].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[0][3].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[0][3].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[0][3].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[0][3].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[0][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[0][3].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[0][4].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[0][4].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[0][4].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[0][4].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[0][4].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[0][4].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[0][4].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[0][4].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[0][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[0][4].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[0][5].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[0][5].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[0][5].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[0][5].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[0][5].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[0][5].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[0][5].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[0][5].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[0][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[0][5].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[0][6].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[0][6].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[0][6].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[0][6].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[0][6].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[0][6].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[0][6].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[0][6].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[0][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[0][6].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[0][7].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[0][7].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[0][7].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[0][7].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[0][7].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[0][7].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[0][7].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[0][7].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[0][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[0][7].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[0][8].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[0][8].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[0][8].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[0][8].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[0][8].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[0][8].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[0][8].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[0][8].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[0][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[0][8].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[0][9].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[0][9].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[0][9].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[0][9].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[0][9].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[0][9].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[0][9].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[0][9].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[0][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[0][9].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[0][10].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[0][10].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[0][10].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[0][10].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[0][10].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[0][10].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[0][10].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[0][10].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[0][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[0][10].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[0][11].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[0][11].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[0][11].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[0][11].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[0][11].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[0][11].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[0][11].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[0][11].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[0][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[0][11].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[0][12].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[0][12].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[0][12].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[0][12].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[0][12].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[0][12].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[0][12].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[0][12].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[0][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[0][12].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[0][13].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[0][13].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[0][13].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[0][13].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[0][13].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[0][13].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[0][13].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[0][13].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[0][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[0][13].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[0][14].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[0][14].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[0][14].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[0][14].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[0][14].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[0][14].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[0][14].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[0][14].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[0][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[0][14].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[0][15].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[0][15].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[0][15].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[0][15].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[0][15].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[0][15].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[0][15].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[0][15].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[0][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[0][15].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[0][16].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[0][16].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[0][16].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[0][16].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[0][16].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[0][16].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[0][16].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[0][16].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[0][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[0][16].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[0][17].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[0][17].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[0][17].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[0][17].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[0][17].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[0][17].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[0][17].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[0][17].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[0][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[0][17].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[0][18].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[0][18].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[0][18].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[0][18].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[0][18].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[0][18].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[0][18].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[0][18].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[0][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[0][18].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[0][19].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[0][19].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[0][19].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[0][19].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[0][19].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[0][19].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[0][19].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[0][19].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[0][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[0][19].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[0][20].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[0][20].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[0][20].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[0][20].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[0][20].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[0][20].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[0][20].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[0][20].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[0][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[0][20].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[0][21].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[0][21].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[0][21].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[0][21].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[0][21].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[0][21].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[0][21].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[0][21].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[0][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[0][21].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[0][22].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[0][22].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[0][22].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[0][22].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[0][22].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[0][22].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[0][22].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[0][22].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[0][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[0][22].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[0][23].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[0][23].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[0][23].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[0][23].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[0][23].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[0][23].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[0][23].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[0][23].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[0][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[0][23].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[0][24].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[0][24].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[0][24].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[0][24].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[0][24].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[0][24].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[0][24].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[0][24].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[0][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[0][24].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[0][25].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[0][25].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[0][25].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[0][25].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[0][25].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[0][25].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[0][25].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[0][25].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[0][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[0][25].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[0][26].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[0][26].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[0][26].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[0][26].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[0][26].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[0][26].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[0][26].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[0][26].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[0][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[0][26].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[0][27].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[0][27].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[0][27].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[0][27].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[0][27].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[0][27].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[0][27].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[0][27].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[0][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[0][27].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[0][28].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[0][28].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[0][28].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[0][28].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[0][28].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[0][28].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[0][28].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[0][28].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[0][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[0][28].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[0][29].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[0][29].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[0][29].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[0][29].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[0][29].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[0][29].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[0][29].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[0][29].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[0][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[0][29].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[0][30].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[0][30].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[0][30].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[0][30].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[0][30].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[0][30].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[0][30].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[0][30].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[0][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[0][30].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[0][31].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[0][31].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[0][31].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[0][31].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[0][31].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[0][31].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[0][31].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[0][31].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[0][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[0][31].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 1
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[1][0].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[1][0].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[1][0].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[1][0].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[1][0].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[1][0].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[1][0].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[1][0].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[1][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[1][0].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[1][1].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[1][1].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[1][1].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[1][1].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[1][1].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[1][1].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[1][1].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[1][1].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[1][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[1][1].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[1][2].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[1][2].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[1][2].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[1][2].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[1][2].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[1][2].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[1][2].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[1][2].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[1][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[1][2].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[1][3].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[1][3].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[1][3].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[1][3].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[1][3].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[1][3].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[1][3].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[1][3].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[1][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[1][3].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[1][4].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[1][4].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[1][4].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[1][4].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[1][4].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[1][4].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[1][4].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[1][4].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[1][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[1][4].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[1][5].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[1][5].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[1][5].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[1][5].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[1][5].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[1][5].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[1][5].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[1][5].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[1][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[1][5].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[1][6].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[1][6].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[1][6].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[1][6].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[1][6].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[1][6].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[1][6].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[1][6].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[1][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[1][6].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[1][7].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[1][7].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[1][7].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[1][7].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[1][7].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[1][7].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[1][7].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[1][7].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[1][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[1][7].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[1][8].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[1][8].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[1][8].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[1][8].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[1][8].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[1][8].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[1][8].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[1][8].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[1][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[1][8].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[1][9].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[1][9].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[1][9].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[1][9].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[1][9].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[1][9].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[1][9].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[1][9].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[1][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[1][9].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[1][10].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[1][10].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[1][10].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[1][10].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[1][10].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[1][10].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[1][10].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[1][10].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[1][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[1][10].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[1][11].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[1][11].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[1][11].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[1][11].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[1][11].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[1][11].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[1][11].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[1][11].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[1][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[1][11].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[1][12].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[1][12].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[1][12].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[1][12].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[1][12].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[1][12].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[1][12].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[1][12].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[1][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[1][12].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[1][13].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[1][13].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[1][13].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[1][13].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[1][13].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[1][13].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[1][13].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[1][13].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[1][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[1][13].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[1][14].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[1][14].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[1][14].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[1][14].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[1][14].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[1][14].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[1][14].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[1][14].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[1][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[1][14].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[1][15].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[1][15].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[1][15].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[1][15].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[1][15].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[1][15].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[1][15].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[1][15].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[1][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[1][15].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[1][16].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[1][16].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[1][16].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[1][16].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[1][16].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[1][16].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[1][16].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[1][16].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[1][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[1][16].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[1][17].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[1][17].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[1][17].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[1][17].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[1][17].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[1][17].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[1][17].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[1][17].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[1][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[1][17].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[1][18].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[1][18].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[1][18].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[1][18].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[1][18].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[1][18].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[1][18].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[1][18].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[1][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[1][18].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[1][19].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[1][19].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[1][19].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[1][19].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[1][19].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[1][19].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[1][19].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[1][19].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[1][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[1][19].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[1][20].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[1][20].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[1][20].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[1][20].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[1][20].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[1][20].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[1][20].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[1][20].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[1][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[1][20].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[1][21].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[1][21].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[1][21].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[1][21].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[1][21].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[1][21].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[1][21].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[1][21].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[1][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[1][21].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[1][22].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[1][22].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[1][22].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[1][22].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[1][22].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[1][22].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[1][22].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[1][22].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[1][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[1][22].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[1][23].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[1][23].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[1][23].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[1][23].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[1][23].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[1][23].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[1][23].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[1][23].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[1][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[1][23].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[1][24].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[1][24].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[1][24].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[1][24].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[1][24].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[1][24].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[1][24].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[1][24].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[1][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[1][24].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[1][25].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[1][25].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[1][25].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[1][25].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[1][25].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[1][25].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[1][25].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[1][25].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[1][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[1][25].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[1][26].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[1][26].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[1][26].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[1][26].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[1][26].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[1][26].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[1][26].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[1][26].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[1][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[1][26].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[1][27].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[1][27].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[1][27].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[1][27].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[1][27].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[1][27].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[1][27].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[1][27].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[1][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[1][27].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[1][28].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[1][28].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[1][28].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[1][28].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[1][28].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[1][28].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[1][28].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[1][28].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[1][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[1][28].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[1][29].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[1][29].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[1][29].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[1][29].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[1][29].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[1][29].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[1][29].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[1][29].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[1][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[1][29].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[1][30].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[1][30].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[1][30].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[1][30].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[1][30].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[1][30].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[1][30].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[1][30].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[1][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[1][30].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[1][31].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[1][31].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[1][31].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[1][31].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[1][31].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[1][31].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[1][31].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[1][31].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[1][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[1][31].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 2
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[2][0].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[2][0].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[2][0].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[2][0].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[2][0].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[2][0].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[2][0].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[2][0].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[2][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[2][0].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[2][1].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[2][1].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[2][1].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[2][1].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[2][1].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[2][1].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[2][1].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[2][1].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[2][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[2][1].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[2][2].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[2][2].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[2][2].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[2][2].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[2][2].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[2][2].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[2][2].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[2][2].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[2][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[2][2].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[2][3].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[2][3].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[2][3].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[2][3].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[2][3].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[2][3].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[2][3].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[2][3].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[2][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[2][3].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[2][4].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[2][4].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[2][4].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[2][4].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[2][4].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[2][4].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[2][4].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[2][4].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[2][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[2][4].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[2][5].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[2][5].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[2][5].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[2][5].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[2][5].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[2][5].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[2][5].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[2][5].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[2][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[2][5].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[2][6].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[2][6].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[2][6].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[2][6].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[2][6].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[2][6].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[2][6].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[2][6].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[2][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[2][6].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[2][7].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[2][7].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[2][7].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[2][7].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[2][7].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[2][7].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[2][7].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[2][7].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[2][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[2][7].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[2][8].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[2][8].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[2][8].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[2][8].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[2][8].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[2][8].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[2][8].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[2][8].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[2][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[2][8].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[2][9].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[2][9].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[2][9].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[2][9].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[2][9].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[2][9].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[2][9].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[2][9].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[2][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[2][9].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[2][10].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[2][10].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[2][10].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[2][10].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[2][10].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[2][10].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[2][10].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[2][10].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[2][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[2][10].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[2][11].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[2][11].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[2][11].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[2][11].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[2][11].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[2][11].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[2][11].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[2][11].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[2][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[2][11].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[2][12].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[2][12].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[2][12].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[2][12].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[2][12].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[2][12].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[2][12].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[2][12].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[2][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[2][12].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[2][13].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[2][13].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[2][13].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[2][13].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[2][13].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[2][13].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[2][13].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[2][13].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[2][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[2][13].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[2][14].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[2][14].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[2][14].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[2][14].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[2][14].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[2][14].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[2][14].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[2][14].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[2][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[2][14].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[2][15].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[2][15].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[2][15].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[2][15].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[2][15].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[2][15].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[2][15].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[2][15].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[2][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[2][15].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[2][16].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[2][16].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[2][16].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[2][16].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[2][16].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[2][16].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[2][16].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[2][16].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[2][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[2][16].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[2][17].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[2][17].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[2][17].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[2][17].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[2][17].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[2][17].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[2][17].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[2][17].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[2][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[2][17].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[2][18].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[2][18].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[2][18].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[2][18].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[2][18].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[2][18].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[2][18].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[2][18].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[2][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[2][18].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[2][19].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[2][19].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[2][19].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[2][19].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[2][19].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[2][19].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[2][19].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[2][19].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[2][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[2][19].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[2][20].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[2][20].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[2][20].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[2][20].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[2][20].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[2][20].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[2][20].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[2][20].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[2][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[2][20].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[2][21].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[2][21].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[2][21].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[2][21].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[2][21].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[2][21].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[2][21].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[2][21].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[2][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[2][21].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[2][22].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[2][22].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[2][22].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[2][22].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[2][22].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[2][22].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[2][22].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[2][22].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[2][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[2][22].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[2][23].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[2][23].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[2][23].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[2][23].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[2][23].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[2][23].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[2][23].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[2][23].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[2][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[2][23].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[2][24].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[2][24].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[2][24].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[2][24].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[2][24].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[2][24].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[2][24].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[2][24].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[2][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[2][24].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[2][25].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[2][25].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[2][25].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[2][25].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[2][25].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[2][25].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[2][25].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[2][25].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[2][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[2][25].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[2][26].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[2][26].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[2][26].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[2][26].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[2][26].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[2][26].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[2][26].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[2][26].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[2][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[2][26].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[2][27].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[2][27].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[2][27].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[2][27].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[2][27].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[2][27].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[2][27].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[2][27].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[2][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[2][27].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[2][28].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[2][28].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[2][28].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[2][28].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[2][28].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[2][28].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[2][28].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[2][28].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[2][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[2][28].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[2][29].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[2][29].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[2][29].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[2][29].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[2][29].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[2][29].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[2][29].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[2][29].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[2][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[2][29].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[2][30].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[2][30].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[2][30].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[2][30].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[2][30].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[2][30].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[2][30].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[2][30].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[2][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[2][30].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[2][31].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[2][31].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[2][31].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[2][31].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[2][31].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[2][31].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[2][31].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[2][31].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[2][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[2][31].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 3
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[3][0].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[3][0].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[3][0].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[3][0].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[3][0].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[3][0].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[3][0].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[3][0].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[3][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[3][0].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[3][1].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[3][1].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[3][1].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[3][1].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[3][1].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[3][1].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[3][1].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[3][1].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[3][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[3][1].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[3][2].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[3][2].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[3][2].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[3][2].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[3][2].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[3][2].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[3][2].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[3][2].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[3][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[3][2].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[3][3].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[3][3].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[3][3].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[3][3].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[3][3].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[3][3].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[3][3].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[3][3].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[3][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[3][3].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[3][4].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[3][4].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[3][4].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[3][4].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[3][4].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[3][4].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[3][4].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[3][4].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[3][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[3][4].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[3][5].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[3][5].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[3][5].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[3][5].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[3][5].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[3][5].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[3][5].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[3][5].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[3][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[3][5].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[3][6].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[3][6].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[3][6].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[3][6].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[3][6].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[3][6].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[3][6].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[3][6].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[3][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[3][6].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[3][7].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[3][7].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[3][7].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[3][7].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[3][7].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[3][7].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[3][7].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[3][7].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[3][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[3][7].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[3][8].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[3][8].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[3][8].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[3][8].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[3][8].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[3][8].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[3][8].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[3][8].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[3][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[3][8].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[3][9].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[3][9].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[3][9].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[3][9].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[3][9].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[3][9].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[3][9].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[3][9].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[3][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[3][9].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[3][10].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[3][10].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[3][10].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[3][10].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[3][10].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[3][10].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[3][10].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[3][10].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[3][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[3][10].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[3][11].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[3][11].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[3][11].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[3][11].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[3][11].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[3][11].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[3][11].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[3][11].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[3][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[3][11].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[3][12].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[3][12].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[3][12].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[3][12].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[3][12].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[3][12].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[3][12].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[3][12].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[3][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[3][12].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[3][13].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[3][13].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[3][13].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[3][13].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[3][13].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[3][13].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[3][13].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[3][13].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[3][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[3][13].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[3][14].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[3][14].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[3][14].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[3][14].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[3][14].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[3][14].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[3][14].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[3][14].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[3][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[3][14].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[3][15].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[3][15].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[3][15].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[3][15].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[3][15].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[3][15].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[3][15].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[3][15].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[3][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[3][15].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[3][16].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[3][16].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[3][16].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[3][16].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[3][16].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[3][16].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[3][16].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[3][16].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[3][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[3][16].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[3][17].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[3][17].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[3][17].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[3][17].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[3][17].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[3][17].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[3][17].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[3][17].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[3][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[3][17].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[3][18].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[3][18].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[3][18].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[3][18].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[3][18].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[3][18].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[3][18].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[3][18].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[3][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[3][18].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[3][19].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[3][19].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[3][19].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[3][19].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[3][19].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[3][19].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[3][19].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[3][19].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[3][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[3][19].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[3][20].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[3][20].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[3][20].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[3][20].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[3][20].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[3][20].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[3][20].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[3][20].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[3][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[3][20].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[3][21].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[3][21].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[3][21].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[3][21].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[3][21].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[3][21].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[3][21].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[3][21].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[3][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[3][21].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[3][22].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[3][22].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[3][22].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[3][22].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[3][22].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[3][22].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[3][22].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[3][22].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[3][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[3][22].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[3][23].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[3][23].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[3][23].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[3][23].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[3][23].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[3][23].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[3][23].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[3][23].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[3][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[3][23].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[3][24].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[3][24].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[3][24].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[3][24].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[3][24].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[3][24].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[3][24].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[3][24].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[3][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[3][24].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[3][25].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[3][25].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[3][25].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[3][25].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[3][25].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[3][25].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[3][25].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[3][25].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[3][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[3][25].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[3][26].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[3][26].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[3][26].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[3][26].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[3][26].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[3][26].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[3][26].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[3][26].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[3][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[3][26].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[3][27].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[3][27].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[3][27].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[3][27].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[3][27].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[3][27].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[3][27].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[3][27].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[3][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[3][27].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[3][28].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[3][28].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[3][28].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[3][28].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[3][28].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[3][28].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[3][28].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[3][28].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[3][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[3][28].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[3][29].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[3][29].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[3][29].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[3][29].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[3][29].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[3][29].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[3][29].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[3][29].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[3][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[3][29].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[3][30].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[3][30].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[3][30].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[3][30].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[3][30].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[3][30].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[3][30].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[3][30].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[3][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[3][30].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[3][31].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[3][31].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[3][31].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[3][31].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[3][31].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[3][31].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[3][31].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[3][31].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[3][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[3][31].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 4
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[4][0].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[4][0].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[4][0].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[4][0].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[4][0].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[4][0].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[4][0].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[4][0].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[4][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[4][0].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[4][1].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[4][1].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[4][1].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[4][1].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[4][1].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[4][1].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[4][1].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[4][1].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[4][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[4][1].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[4][2].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[4][2].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[4][2].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[4][2].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[4][2].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[4][2].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[4][2].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[4][2].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[4][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[4][2].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[4][3].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[4][3].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[4][3].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[4][3].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[4][3].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[4][3].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[4][3].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[4][3].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[4][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[4][3].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[4][4].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[4][4].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[4][4].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[4][4].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[4][4].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[4][4].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[4][4].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[4][4].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[4][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[4][4].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[4][5].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[4][5].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[4][5].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[4][5].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[4][5].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[4][5].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[4][5].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[4][5].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[4][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[4][5].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[4][6].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[4][6].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[4][6].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[4][6].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[4][6].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[4][6].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[4][6].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[4][6].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[4][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[4][6].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[4][7].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[4][7].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[4][7].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[4][7].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[4][7].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[4][7].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[4][7].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[4][7].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[4][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[4][7].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[4][8].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[4][8].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[4][8].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[4][8].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[4][8].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[4][8].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[4][8].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[4][8].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[4][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[4][8].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[4][9].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[4][9].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[4][9].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[4][9].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[4][9].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[4][9].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[4][9].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[4][9].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[4][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[4][9].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[4][10].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[4][10].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[4][10].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[4][10].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[4][10].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[4][10].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[4][10].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[4][10].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[4][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[4][10].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[4][11].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[4][11].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[4][11].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[4][11].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[4][11].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[4][11].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[4][11].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[4][11].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[4][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[4][11].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[4][12].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[4][12].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[4][12].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[4][12].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[4][12].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[4][12].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[4][12].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[4][12].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[4][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[4][12].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[4][13].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[4][13].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[4][13].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[4][13].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[4][13].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[4][13].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[4][13].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[4][13].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[4][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[4][13].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[4][14].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[4][14].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[4][14].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[4][14].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[4][14].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[4][14].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[4][14].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[4][14].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[4][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[4][14].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[4][15].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[4][15].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[4][15].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[4][15].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[4][15].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[4][15].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[4][15].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[4][15].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[4][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[4][15].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[4][16].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[4][16].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[4][16].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[4][16].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[4][16].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[4][16].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[4][16].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[4][16].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[4][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[4][16].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[4][17].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[4][17].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[4][17].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[4][17].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[4][17].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[4][17].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[4][17].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[4][17].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[4][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[4][17].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[4][18].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[4][18].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[4][18].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[4][18].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[4][18].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[4][18].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[4][18].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[4][18].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[4][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[4][18].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[4][19].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[4][19].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[4][19].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[4][19].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[4][19].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[4][19].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[4][19].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[4][19].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[4][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[4][19].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[4][20].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[4][20].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[4][20].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[4][20].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[4][20].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[4][20].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[4][20].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[4][20].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[4][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[4][20].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[4][21].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[4][21].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[4][21].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[4][21].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[4][21].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[4][21].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[4][21].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[4][21].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[4][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[4][21].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[4][22].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[4][22].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[4][22].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[4][22].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[4][22].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[4][22].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[4][22].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[4][22].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[4][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[4][22].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[4][23].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[4][23].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[4][23].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[4][23].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[4][23].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[4][23].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[4][23].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[4][23].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[4][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[4][23].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[4][24].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[4][24].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[4][24].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[4][24].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[4][24].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[4][24].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[4][24].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[4][24].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[4][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[4][24].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[4][25].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[4][25].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[4][25].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[4][25].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[4][25].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[4][25].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[4][25].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[4][25].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[4][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[4][25].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[4][26].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[4][26].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[4][26].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[4][26].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[4][26].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[4][26].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[4][26].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[4][26].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[4][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[4][26].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[4][27].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[4][27].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[4][27].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[4][27].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[4][27].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[4][27].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[4][27].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[4][27].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[4][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[4][27].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[4][28].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[4][28].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[4][28].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[4][28].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[4][28].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[4][28].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[4][28].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[4][28].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[4][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[4][28].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[4][29].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[4][29].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[4][29].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[4][29].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[4][29].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[4][29].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[4][29].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[4][29].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[4][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[4][29].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[4][30].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[4][30].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[4][30].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[4][30].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[4][30].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[4][30].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[4][30].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[4][30].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[4][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[4][30].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[4][31].dma__memc__write_valid      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[4][31].dma__memc__write_address    = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[4][31].dma__memc__write_data       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[4][31].dma__memc__read_valid       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[4][31].dma__memc__read_address     = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[4][31].dma__memc__read_pause       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[4][31].memc__dma__write_ready      = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[4][31].memc__dma__read_data        = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[4][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[4][31].memc__dma__read_ready       = pe_array_inst.pe_inst[4].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 5
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[5][0].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[5][0].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[5][0].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[5][0].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[5][0].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[5][0].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[5][0].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[5][0].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[5][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[5][0].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[5][1].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[5][1].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[5][1].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[5][1].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[5][1].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[5][1].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[5][1].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[5][1].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[5][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[5][1].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[5][2].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[5][2].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[5][2].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[5][2].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[5][2].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[5][2].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[5][2].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[5][2].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[5][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[5][2].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[5][3].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[5][3].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[5][3].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[5][3].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[5][3].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[5][3].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[5][3].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[5][3].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[5][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[5][3].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[5][4].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[5][4].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[5][4].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[5][4].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[5][4].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[5][4].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[5][4].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[5][4].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[5][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[5][4].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[5][5].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[5][5].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[5][5].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[5][5].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[5][5].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[5][5].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[5][5].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[5][5].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[5][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[5][5].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[5][6].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[5][6].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[5][6].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[5][6].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[5][6].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[5][6].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[5][6].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[5][6].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[5][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[5][6].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[5][7].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[5][7].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[5][7].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[5][7].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[5][7].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[5][7].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[5][7].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[5][7].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[5][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[5][7].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[5][8].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[5][8].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[5][8].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[5][8].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[5][8].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[5][8].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[5][8].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[5][8].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[5][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[5][8].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[5][9].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[5][9].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[5][9].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[5][9].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[5][9].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[5][9].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[5][9].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[5][9].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[5][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[5][9].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[5][10].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[5][10].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[5][10].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[5][10].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[5][10].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[5][10].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[5][10].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[5][10].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[5][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[5][10].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[5][11].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[5][11].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[5][11].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[5][11].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[5][11].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[5][11].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[5][11].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[5][11].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[5][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[5][11].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[5][12].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[5][12].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[5][12].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[5][12].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[5][12].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[5][12].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[5][12].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[5][12].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[5][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[5][12].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[5][13].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[5][13].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[5][13].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[5][13].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[5][13].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[5][13].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[5][13].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[5][13].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[5][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[5][13].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[5][14].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[5][14].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[5][14].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[5][14].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[5][14].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[5][14].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[5][14].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[5][14].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[5][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[5][14].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[5][15].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[5][15].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[5][15].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[5][15].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[5][15].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[5][15].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[5][15].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[5][15].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[5][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[5][15].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[5][16].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[5][16].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[5][16].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[5][16].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[5][16].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[5][16].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[5][16].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[5][16].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[5][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[5][16].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[5][17].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[5][17].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[5][17].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[5][17].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[5][17].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[5][17].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[5][17].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[5][17].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[5][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[5][17].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[5][18].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[5][18].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[5][18].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[5][18].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[5][18].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[5][18].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[5][18].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[5][18].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[5][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[5][18].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[5][19].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[5][19].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[5][19].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[5][19].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[5][19].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[5][19].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[5][19].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[5][19].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[5][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[5][19].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[5][20].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[5][20].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[5][20].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[5][20].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[5][20].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[5][20].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[5][20].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[5][20].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[5][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[5][20].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[5][21].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[5][21].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[5][21].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[5][21].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[5][21].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[5][21].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[5][21].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[5][21].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[5][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[5][21].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[5][22].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[5][22].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[5][22].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[5][22].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[5][22].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[5][22].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[5][22].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[5][22].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[5][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[5][22].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[5][23].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[5][23].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[5][23].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[5][23].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[5][23].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[5][23].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[5][23].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[5][23].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[5][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[5][23].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[5][24].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[5][24].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[5][24].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[5][24].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[5][24].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[5][24].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[5][24].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[5][24].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[5][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[5][24].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[5][25].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[5][25].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[5][25].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[5][25].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[5][25].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[5][25].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[5][25].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[5][25].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[5][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[5][25].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[5][26].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[5][26].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[5][26].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[5][26].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[5][26].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[5][26].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[5][26].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[5][26].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[5][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[5][26].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[5][27].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[5][27].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[5][27].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[5][27].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[5][27].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[5][27].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[5][27].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[5][27].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[5][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[5][27].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[5][28].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[5][28].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[5][28].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[5][28].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[5][28].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[5][28].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[5][28].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[5][28].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[5][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[5][28].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[5][29].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[5][29].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[5][29].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[5][29].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[5][29].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[5][29].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[5][29].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[5][29].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[5][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[5][29].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[5][30].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[5][30].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[5][30].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[5][30].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[5][30].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[5][30].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[5][30].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[5][30].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[5][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[5][30].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[5][31].dma__memc__write_valid      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[5][31].dma__memc__write_address    = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[5][31].dma__memc__write_data       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[5][31].dma__memc__read_valid       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[5][31].dma__memc__read_address     = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[5][31].dma__memc__read_pause       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[5][31].memc__dma__write_ready      = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[5][31].memc__dma__read_data        = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[5][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[5][31].memc__dma__read_ready       = pe_array_inst.pe_inst[5].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 6
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[6][0].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[6][0].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[6][0].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[6][0].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[6][0].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[6][0].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[6][0].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[6][0].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[6][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[6][0].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[6][1].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[6][1].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[6][1].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[6][1].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[6][1].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[6][1].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[6][1].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[6][1].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[6][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[6][1].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[6][2].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[6][2].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[6][2].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[6][2].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[6][2].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[6][2].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[6][2].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[6][2].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[6][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[6][2].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[6][3].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[6][3].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[6][3].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[6][3].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[6][3].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[6][3].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[6][3].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[6][3].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[6][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[6][3].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[6][4].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[6][4].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[6][4].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[6][4].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[6][4].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[6][4].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[6][4].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[6][4].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[6][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[6][4].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[6][5].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[6][5].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[6][5].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[6][5].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[6][5].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[6][5].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[6][5].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[6][5].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[6][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[6][5].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[6][6].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[6][6].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[6][6].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[6][6].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[6][6].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[6][6].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[6][6].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[6][6].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[6][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[6][6].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[6][7].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[6][7].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[6][7].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[6][7].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[6][7].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[6][7].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[6][7].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[6][7].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[6][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[6][7].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[6][8].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[6][8].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[6][8].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[6][8].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[6][8].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[6][8].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[6][8].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[6][8].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[6][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[6][8].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[6][9].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[6][9].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[6][9].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[6][9].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[6][9].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[6][9].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[6][9].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[6][9].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[6][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[6][9].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[6][10].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[6][10].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[6][10].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[6][10].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[6][10].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[6][10].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[6][10].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[6][10].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[6][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[6][10].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[6][11].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[6][11].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[6][11].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[6][11].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[6][11].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[6][11].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[6][11].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[6][11].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[6][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[6][11].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[6][12].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[6][12].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[6][12].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[6][12].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[6][12].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[6][12].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[6][12].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[6][12].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[6][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[6][12].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[6][13].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[6][13].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[6][13].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[6][13].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[6][13].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[6][13].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[6][13].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[6][13].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[6][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[6][13].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[6][14].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[6][14].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[6][14].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[6][14].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[6][14].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[6][14].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[6][14].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[6][14].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[6][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[6][14].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[6][15].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[6][15].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[6][15].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[6][15].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[6][15].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[6][15].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[6][15].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[6][15].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[6][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[6][15].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[6][16].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[6][16].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[6][16].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[6][16].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[6][16].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[6][16].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[6][16].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[6][16].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[6][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[6][16].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[6][17].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[6][17].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[6][17].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[6][17].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[6][17].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[6][17].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[6][17].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[6][17].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[6][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[6][17].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[6][18].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[6][18].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[6][18].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[6][18].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[6][18].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[6][18].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[6][18].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[6][18].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[6][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[6][18].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[6][19].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[6][19].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[6][19].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[6][19].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[6][19].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[6][19].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[6][19].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[6][19].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[6][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[6][19].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[6][20].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[6][20].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[6][20].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[6][20].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[6][20].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[6][20].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[6][20].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[6][20].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[6][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[6][20].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[6][21].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[6][21].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[6][21].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[6][21].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[6][21].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[6][21].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[6][21].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[6][21].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[6][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[6][21].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[6][22].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[6][22].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[6][22].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[6][22].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[6][22].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[6][22].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[6][22].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[6][22].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[6][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[6][22].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[6][23].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[6][23].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[6][23].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[6][23].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[6][23].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[6][23].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[6][23].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[6][23].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[6][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[6][23].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[6][24].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[6][24].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[6][24].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[6][24].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[6][24].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[6][24].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[6][24].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[6][24].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[6][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[6][24].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[6][25].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[6][25].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[6][25].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[6][25].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[6][25].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[6][25].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[6][25].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[6][25].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[6][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[6][25].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[6][26].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[6][26].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[6][26].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[6][26].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[6][26].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[6][26].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[6][26].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[6][26].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[6][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[6][26].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[6][27].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[6][27].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[6][27].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[6][27].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[6][27].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[6][27].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[6][27].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[6][27].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[6][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[6][27].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[6][28].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[6][28].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[6][28].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[6][28].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[6][28].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[6][28].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[6][28].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[6][28].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[6][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[6][28].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[6][29].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[6][29].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[6][29].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[6][29].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[6][29].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[6][29].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[6][29].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[6][29].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[6][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[6][29].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[6][30].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[6][30].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[6][30].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[6][30].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[6][30].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[6][30].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[6][30].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[6][30].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[6][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[6][30].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[6][31].dma__memc__write_valid      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[6][31].dma__memc__write_address    = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[6][31].dma__memc__write_data       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[6][31].dma__memc__read_valid       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[6][31].dma__memc__read_address     = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[6][31].dma__memc__read_pause       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[6][31].memc__dma__write_ready      = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[6][31].memc__dma__read_data        = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[6][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[6][31].memc__dma__read_ready       = pe_array_inst.pe_inst[6].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 7
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[7][0].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[7][0].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[7][0].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[7][0].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[7][0].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[7][0].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[7][0].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[7][0].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[7][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[7][0].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[7][1].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[7][1].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[7][1].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[7][1].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[7][1].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[7][1].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[7][1].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[7][1].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[7][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[7][1].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[7][2].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[7][2].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[7][2].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[7][2].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[7][2].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[7][2].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[7][2].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[7][2].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[7][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[7][2].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[7][3].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[7][3].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[7][3].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[7][3].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[7][3].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[7][3].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[7][3].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[7][3].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[7][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[7][3].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[7][4].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[7][4].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[7][4].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[7][4].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[7][4].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[7][4].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[7][4].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[7][4].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[7][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[7][4].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[7][5].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[7][5].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[7][5].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[7][5].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[7][5].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[7][5].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[7][5].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[7][5].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[7][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[7][5].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[7][6].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[7][6].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[7][6].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[7][6].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[7][6].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[7][6].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[7][6].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[7][6].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[7][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[7][6].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[7][7].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[7][7].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[7][7].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[7][7].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[7][7].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[7][7].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[7][7].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[7][7].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[7][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[7][7].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[7][8].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[7][8].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[7][8].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[7][8].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[7][8].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[7][8].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[7][8].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[7][8].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[7][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[7][8].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[7][9].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[7][9].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[7][9].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[7][9].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[7][9].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[7][9].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[7][9].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[7][9].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[7][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[7][9].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[7][10].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[7][10].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[7][10].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[7][10].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[7][10].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[7][10].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[7][10].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[7][10].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[7][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[7][10].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[7][11].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[7][11].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[7][11].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[7][11].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[7][11].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[7][11].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[7][11].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[7][11].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[7][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[7][11].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[7][12].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[7][12].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[7][12].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[7][12].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[7][12].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[7][12].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[7][12].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[7][12].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[7][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[7][12].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[7][13].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[7][13].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[7][13].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[7][13].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[7][13].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[7][13].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[7][13].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[7][13].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[7][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[7][13].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[7][14].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[7][14].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[7][14].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[7][14].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[7][14].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[7][14].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[7][14].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[7][14].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[7][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[7][14].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[7][15].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[7][15].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[7][15].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[7][15].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[7][15].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[7][15].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[7][15].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[7][15].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[7][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[7][15].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[7][16].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[7][16].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[7][16].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[7][16].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[7][16].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[7][16].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[7][16].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[7][16].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[7][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[7][16].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[7][17].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[7][17].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[7][17].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[7][17].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[7][17].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[7][17].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[7][17].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[7][17].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[7][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[7][17].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[7][18].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[7][18].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[7][18].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[7][18].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[7][18].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[7][18].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[7][18].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[7][18].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[7][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[7][18].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[7][19].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[7][19].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[7][19].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[7][19].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[7][19].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[7][19].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[7][19].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[7][19].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[7][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[7][19].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[7][20].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[7][20].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[7][20].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[7][20].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[7][20].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[7][20].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[7][20].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[7][20].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[7][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[7][20].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[7][21].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[7][21].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[7][21].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[7][21].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[7][21].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[7][21].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[7][21].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[7][21].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[7][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[7][21].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[7][22].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[7][22].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[7][22].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[7][22].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[7][22].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[7][22].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[7][22].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[7][22].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[7][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[7][22].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[7][23].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[7][23].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[7][23].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[7][23].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[7][23].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[7][23].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[7][23].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[7][23].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[7][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[7][23].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[7][24].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[7][24].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[7][24].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[7][24].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[7][24].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[7][24].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[7][24].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[7][24].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[7][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[7][24].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[7][25].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[7][25].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[7][25].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[7][25].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[7][25].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[7][25].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[7][25].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[7][25].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[7][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[7][25].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[7][26].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[7][26].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[7][26].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[7][26].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[7][26].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[7][26].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[7][26].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[7][26].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[7][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[7][26].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[7][27].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[7][27].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[7][27].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[7][27].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[7][27].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[7][27].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[7][27].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[7][27].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[7][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[7][27].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[7][28].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[7][28].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[7][28].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[7][28].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[7][28].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[7][28].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[7][28].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[7][28].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[7][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[7][28].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[7][29].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[7][29].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[7][29].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[7][29].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[7][29].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[7][29].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[7][29].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[7][29].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[7][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[7][29].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[7][30].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[7][30].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[7][30].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[7][30].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[7][30].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[7][30].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[7][30].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[7][30].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[7][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[7][30].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[7][31].dma__memc__write_valid      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[7][31].dma__memc__write_address    = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[7][31].dma__memc__write_data       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[7][31].dma__memc__read_valid       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[7][31].dma__memc__read_address     = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[7][31].dma__memc__read_pause       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[7][31].memc__dma__write_ready      = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[7][31].memc__dma__read_data        = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[7][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[7][31].memc__dma__read_ready       = pe_array_inst.pe_inst[7].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 8
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[8][0].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[8][0].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[8][0].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[8][0].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[8][0].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[8][0].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[8][0].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[8][0].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[8][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[8][0].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[8][1].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[8][1].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[8][1].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[8][1].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[8][1].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[8][1].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[8][1].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[8][1].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[8][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[8][1].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[8][2].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[8][2].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[8][2].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[8][2].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[8][2].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[8][2].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[8][2].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[8][2].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[8][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[8][2].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[8][3].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[8][3].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[8][3].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[8][3].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[8][3].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[8][3].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[8][3].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[8][3].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[8][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[8][3].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[8][4].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[8][4].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[8][4].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[8][4].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[8][4].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[8][4].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[8][4].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[8][4].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[8][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[8][4].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[8][5].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[8][5].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[8][5].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[8][5].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[8][5].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[8][5].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[8][5].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[8][5].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[8][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[8][5].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[8][6].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[8][6].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[8][6].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[8][6].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[8][6].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[8][6].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[8][6].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[8][6].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[8][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[8][6].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[8][7].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[8][7].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[8][7].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[8][7].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[8][7].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[8][7].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[8][7].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[8][7].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[8][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[8][7].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[8][8].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[8][8].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[8][8].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[8][8].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[8][8].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[8][8].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[8][8].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[8][8].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[8][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[8][8].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[8][9].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[8][9].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[8][9].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[8][9].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[8][9].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[8][9].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[8][9].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[8][9].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[8][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[8][9].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[8][10].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[8][10].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[8][10].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[8][10].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[8][10].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[8][10].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[8][10].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[8][10].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[8][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[8][10].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[8][11].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[8][11].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[8][11].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[8][11].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[8][11].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[8][11].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[8][11].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[8][11].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[8][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[8][11].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[8][12].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[8][12].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[8][12].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[8][12].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[8][12].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[8][12].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[8][12].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[8][12].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[8][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[8][12].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[8][13].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[8][13].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[8][13].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[8][13].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[8][13].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[8][13].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[8][13].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[8][13].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[8][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[8][13].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[8][14].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[8][14].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[8][14].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[8][14].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[8][14].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[8][14].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[8][14].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[8][14].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[8][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[8][14].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[8][15].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[8][15].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[8][15].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[8][15].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[8][15].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[8][15].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[8][15].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[8][15].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[8][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[8][15].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[8][16].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[8][16].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[8][16].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[8][16].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[8][16].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[8][16].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[8][16].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[8][16].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[8][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[8][16].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[8][17].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[8][17].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[8][17].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[8][17].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[8][17].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[8][17].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[8][17].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[8][17].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[8][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[8][17].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[8][18].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[8][18].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[8][18].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[8][18].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[8][18].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[8][18].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[8][18].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[8][18].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[8][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[8][18].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[8][19].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[8][19].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[8][19].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[8][19].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[8][19].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[8][19].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[8][19].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[8][19].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[8][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[8][19].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[8][20].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[8][20].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[8][20].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[8][20].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[8][20].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[8][20].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[8][20].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[8][20].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[8][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[8][20].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[8][21].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[8][21].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[8][21].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[8][21].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[8][21].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[8][21].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[8][21].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[8][21].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[8][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[8][21].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[8][22].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[8][22].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[8][22].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[8][22].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[8][22].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[8][22].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[8][22].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[8][22].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[8][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[8][22].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[8][23].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[8][23].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[8][23].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[8][23].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[8][23].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[8][23].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[8][23].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[8][23].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[8][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[8][23].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[8][24].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[8][24].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[8][24].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[8][24].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[8][24].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[8][24].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[8][24].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[8][24].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[8][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[8][24].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[8][25].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[8][25].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[8][25].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[8][25].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[8][25].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[8][25].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[8][25].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[8][25].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[8][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[8][25].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[8][26].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[8][26].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[8][26].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[8][26].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[8][26].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[8][26].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[8][26].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[8][26].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[8][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[8][26].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[8][27].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[8][27].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[8][27].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[8][27].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[8][27].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[8][27].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[8][27].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[8][27].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[8][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[8][27].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[8][28].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[8][28].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[8][28].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[8][28].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[8][28].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[8][28].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[8][28].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[8][28].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[8][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[8][28].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[8][29].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[8][29].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[8][29].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[8][29].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[8][29].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[8][29].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[8][29].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[8][29].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[8][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[8][29].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[8][30].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[8][30].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[8][30].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[8][30].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[8][30].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[8][30].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[8][30].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[8][30].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[8][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[8][30].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[8][31].dma__memc__write_valid      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[8][31].dma__memc__write_address    = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[8][31].dma__memc__write_data       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[8][31].dma__memc__read_valid       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[8][31].dma__memc__read_address     = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[8][31].dma__memc__read_pause       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[8][31].memc__dma__write_ready      = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[8][31].memc__dma__read_data        = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[8][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[8][31].memc__dma__read_ready       = pe_array_inst.pe_inst[8].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 9
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[9][0].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[9][0].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[9][0].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[9][0].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[9][0].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[9][0].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[9][0].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[9][0].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[9][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[9][0].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[9][1].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[9][1].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[9][1].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[9][1].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[9][1].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[9][1].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[9][1].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[9][1].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[9][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[9][1].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[9][2].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[9][2].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[9][2].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[9][2].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[9][2].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[9][2].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[9][2].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[9][2].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[9][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[9][2].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[9][3].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[9][3].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[9][3].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[9][3].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[9][3].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[9][3].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[9][3].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[9][3].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[9][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[9][3].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[9][4].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[9][4].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[9][4].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[9][4].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[9][4].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[9][4].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[9][4].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[9][4].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[9][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[9][4].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[9][5].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[9][5].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[9][5].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[9][5].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[9][5].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[9][5].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[9][5].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[9][5].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[9][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[9][5].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[9][6].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[9][6].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[9][6].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[9][6].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[9][6].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[9][6].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[9][6].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[9][6].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[9][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[9][6].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[9][7].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[9][7].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[9][7].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[9][7].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[9][7].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[9][7].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[9][7].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[9][7].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[9][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[9][7].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[9][8].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[9][8].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[9][8].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[9][8].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[9][8].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[9][8].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[9][8].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[9][8].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[9][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[9][8].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[9][9].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[9][9].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[9][9].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[9][9].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[9][9].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[9][9].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[9][9].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[9][9].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[9][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[9][9].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[9][10].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[9][10].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[9][10].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[9][10].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[9][10].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[9][10].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[9][10].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[9][10].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[9][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[9][10].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[9][11].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[9][11].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[9][11].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[9][11].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[9][11].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[9][11].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[9][11].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[9][11].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[9][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[9][11].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[9][12].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[9][12].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[9][12].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[9][12].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[9][12].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[9][12].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[9][12].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[9][12].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[9][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[9][12].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[9][13].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[9][13].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[9][13].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[9][13].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[9][13].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[9][13].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[9][13].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[9][13].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[9][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[9][13].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[9][14].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[9][14].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[9][14].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[9][14].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[9][14].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[9][14].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[9][14].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[9][14].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[9][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[9][14].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[9][15].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[9][15].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[9][15].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[9][15].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[9][15].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[9][15].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[9][15].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[9][15].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[9][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[9][15].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[9][16].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[9][16].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[9][16].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[9][16].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[9][16].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[9][16].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[9][16].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[9][16].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[9][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[9][16].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[9][17].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[9][17].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[9][17].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[9][17].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[9][17].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[9][17].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[9][17].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[9][17].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[9][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[9][17].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[9][18].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[9][18].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[9][18].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[9][18].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[9][18].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[9][18].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[9][18].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[9][18].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[9][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[9][18].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[9][19].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[9][19].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[9][19].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[9][19].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[9][19].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[9][19].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[9][19].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[9][19].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[9][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[9][19].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[9][20].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[9][20].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[9][20].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[9][20].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[9][20].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[9][20].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[9][20].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[9][20].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[9][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[9][20].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[9][21].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[9][21].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[9][21].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[9][21].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[9][21].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[9][21].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[9][21].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[9][21].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[9][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[9][21].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[9][22].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[9][22].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[9][22].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[9][22].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[9][22].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[9][22].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[9][22].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[9][22].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[9][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[9][22].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[9][23].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[9][23].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[9][23].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[9][23].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[9][23].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[9][23].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[9][23].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[9][23].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[9][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[9][23].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[9][24].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[9][24].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[9][24].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[9][24].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[9][24].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[9][24].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[9][24].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[9][24].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[9][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[9][24].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[9][25].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[9][25].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[9][25].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[9][25].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[9][25].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[9][25].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[9][25].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[9][25].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[9][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[9][25].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[9][26].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[9][26].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[9][26].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[9][26].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[9][26].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[9][26].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[9][26].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[9][26].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[9][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[9][26].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[9][27].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[9][27].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[9][27].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[9][27].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[9][27].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[9][27].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[9][27].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[9][27].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[9][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[9][27].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[9][28].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[9][28].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[9][28].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[9][28].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[9][28].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[9][28].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[9][28].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[9][28].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[9][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[9][28].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[9][29].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[9][29].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[9][29].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[9][29].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[9][29].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[9][29].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[9][29].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[9][29].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[9][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[9][29].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[9][30].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[9][30].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[9][30].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[9][30].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[9][30].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[9][30].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[9][30].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[9][30].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[9][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[9][30].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[9][31].dma__memc__write_valid      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[9][31].dma__memc__write_address    = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[9][31].dma__memc__write_data       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[9][31].dma__memc__read_valid       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[9][31].dma__memc__read_address     = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[9][31].dma__memc__read_pause       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[9][31].memc__dma__write_ready      = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[9][31].memc__dma__read_data        = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[9][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[9][31].memc__dma__read_ready       = pe_array_inst.pe_inst[9].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 10
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[10][0].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[10][0].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[10][0].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[10][0].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[10][0].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[10][0].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[10][0].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[10][0].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[10][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[10][0].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[10][1].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[10][1].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[10][1].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[10][1].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[10][1].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[10][1].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[10][1].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[10][1].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[10][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[10][1].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[10][2].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[10][2].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[10][2].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[10][2].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[10][2].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[10][2].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[10][2].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[10][2].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[10][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[10][2].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[10][3].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[10][3].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[10][3].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[10][3].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[10][3].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[10][3].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[10][3].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[10][3].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[10][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[10][3].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[10][4].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[10][4].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[10][4].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[10][4].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[10][4].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[10][4].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[10][4].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[10][4].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[10][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[10][4].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[10][5].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[10][5].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[10][5].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[10][5].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[10][5].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[10][5].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[10][5].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[10][5].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[10][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[10][5].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[10][6].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[10][6].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[10][6].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[10][6].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[10][6].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[10][6].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[10][6].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[10][6].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[10][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[10][6].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[10][7].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[10][7].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[10][7].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[10][7].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[10][7].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[10][7].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[10][7].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[10][7].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[10][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[10][7].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[10][8].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[10][8].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[10][8].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[10][8].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[10][8].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[10][8].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[10][8].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[10][8].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[10][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[10][8].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[10][9].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[10][9].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[10][9].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[10][9].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[10][9].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[10][9].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[10][9].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[10][9].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[10][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[10][9].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[10][10].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[10][10].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[10][10].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[10][10].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[10][10].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[10][10].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[10][10].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[10][10].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[10][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[10][10].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[10][11].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[10][11].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[10][11].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[10][11].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[10][11].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[10][11].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[10][11].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[10][11].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[10][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[10][11].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[10][12].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[10][12].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[10][12].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[10][12].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[10][12].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[10][12].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[10][12].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[10][12].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[10][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[10][12].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[10][13].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[10][13].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[10][13].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[10][13].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[10][13].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[10][13].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[10][13].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[10][13].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[10][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[10][13].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[10][14].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[10][14].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[10][14].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[10][14].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[10][14].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[10][14].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[10][14].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[10][14].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[10][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[10][14].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[10][15].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[10][15].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[10][15].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[10][15].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[10][15].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[10][15].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[10][15].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[10][15].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[10][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[10][15].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[10][16].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[10][16].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[10][16].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[10][16].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[10][16].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[10][16].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[10][16].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[10][16].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[10][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[10][16].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[10][17].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[10][17].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[10][17].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[10][17].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[10][17].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[10][17].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[10][17].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[10][17].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[10][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[10][17].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[10][18].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[10][18].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[10][18].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[10][18].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[10][18].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[10][18].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[10][18].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[10][18].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[10][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[10][18].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[10][19].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[10][19].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[10][19].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[10][19].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[10][19].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[10][19].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[10][19].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[10][19].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[10][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[10][19].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[10][20].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[10][20].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[10][20].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[10][20].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[10][20].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[10][20].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[10][20].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[10][20].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[10][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[10][20].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[10][21].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[10][21].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[10][21].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[10][21].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[10][21].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[10][21].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[10][21].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[10][21].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[10][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[10][21].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[10][22].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[10][22].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[10][22].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[10][22].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[10][22].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[10][22].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[10][22].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[10][22].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[10][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[10][22].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[10][23].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[10][23].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[10][23].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[10][23].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[10][23].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[10][23].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[10][23].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[10][23].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[10][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[10][23].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[10][24].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[10][24].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[10][24].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[10][24].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[10][24].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[10][24].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[10][24].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[10][24].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[10][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[10][24].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[10][25].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[10][25].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[10][25].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[10][25].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[10][25].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[10][25].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[10][25].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[10][25].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[10][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[10][25].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[10][26].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[10][26].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[10][26].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[10][26].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[10][26].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[10][26].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[10][26].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[10][26].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[10][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[10][26].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[10][27].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[10][27].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[10][27].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[10][27].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[10][27].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[10][27].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[10][27].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[10][27].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[10][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[10][27].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[10][28].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[10][28].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[10][28].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[10][28].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[10][28].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[10][28].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[10][28].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[10][28].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[10][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[10][28].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[10][29].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[10][29].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[10][29].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[10][29].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[10][29].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[10][29].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[10][29].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[10][29].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[10][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[10][29].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[10][30].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[10][30].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[10][30].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[10][30].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[10][30].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[10][30].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[10][30].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[10][30].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[10][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[10][30].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[10][31].dma__memc__write_valid      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[10][31].dma__memc__write_address    = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[10][31].dma__memc__write_data       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[10][31].dma__memc__read_valid       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[10][31].dma__memc__read_address     = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[10][31].dma__memc__read_pause       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[10][31].memc__dma__write_ready      = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[10][31].memc__dma__read_data        = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[10][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[10][31].memc__dma__read_ready       = pe_array_inst.pe_inst[10].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 11
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[11][0].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[11][0].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[11][0].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[11][0].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[11][0].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[11][0].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[11][0].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[11][0].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[11][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[11][0].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[11][1].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[11][1].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[11][1].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[11][1].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[11][1].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[11][1].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[11][1].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[11][1].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[11][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[11][1].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[11][2].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[11][2].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[11][2].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[11][2].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[11][2].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[11][2].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[11][2].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[11][2].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[11][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[11][2].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[11][3].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[11][3].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[11][3].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[11][3].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[11][3].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[11][3].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[11][3].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[11][3].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[11][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[11][3].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[11][4].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[11][4].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[11][4].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[11][4].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[11][4].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[11][4].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[11][4].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[11][4].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[11][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[11][4].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[11][5].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[11][5].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[11][5].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[11][5].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[11][5].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[11][5].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[11][5].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[11][5].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[11][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[11][5].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[11][6].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[11][6].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[11][6].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[11][6].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[11][6].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[11][6].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[11][6].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[11][6].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[11][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[11][6].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[11][7].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[11][7].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[11][7].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[11][7].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[11][7].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[11][7].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[11][7].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[11][7].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[11][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[11][7].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[11][8].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[11][8].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[11][8].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[11][8].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[11][8].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[11][8].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[11][8].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[11][8].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[11][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[11][8].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[11][9].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[11][9].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[11][9].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[11][9].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[11][9].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[11][9].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[11][9].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[11][9].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[11][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[11][9].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[11][10].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[11][10].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[11][10].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[11][10].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[11][10].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[11][10].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[11][10].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[11][10].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[11][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[11][10].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[11][11].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[11][11].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[11][11].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[11][11].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[11][11].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[11][11].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[11][11].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[11][11].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[11][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[11][11].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[11][12].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[11][12].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[11][12].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[11][12].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[11][12].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[11][12].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[11][12].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[11][12].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[11][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[11][12].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[11][13].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[11][13].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[11][13].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[11][13].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[11][13].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[11][13].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[11][13].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[11][13].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[11][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[11][13].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[11][14].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[11][14].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[11][14].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[11][14].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[11][14].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[11][14].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[11][14].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[11][14].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[11][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[11][14].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[11][15].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[11][15].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[11][15].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[11][15].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[11][15].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[11][15].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[11][15].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[11][15].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[11][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[11][15].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[11][16].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[11][16].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[11][16].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[11][16].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[11][16].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[11][16].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[11][16].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[11][16].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[11][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[11][16].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[11][17].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[11][17].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[11][17].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[11][17].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[11][17].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[11][17].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[11][17].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[11][17].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[11][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[11][17].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[11][18].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[11][18].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[11][18].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[11][18].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[11][18].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[11][18].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[11][18].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[11][18].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[11][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[11][18].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[11][19].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[11][19].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[11][19].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[11][19].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[11][19].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[11][19].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[11][19].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[11][19].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[11][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[11][19].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[11][20].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[11][20].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[11][20].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[11][20].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[11][20].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[11][20].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[11][20].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[11][20].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[11][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[11][20].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[11][21].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[11][21].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[11][21].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[11][21].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[11][21].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[11][21].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[11][21].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[11][21].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[11][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[11][21].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[11][22].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[11][22].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[11][22].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[11][22].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[11][22].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[11][22].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[11][22].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[11][22].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[11][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[11][22].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[11][23].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[11][23].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[11][23].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[11][23].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[11][23].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[11][23].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[11][23].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[11][23].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[11][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[11][23].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[11][24].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[11][24].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[11][24].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[11][24].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[11][24].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[11][24].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[11][24].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[11][24].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[11][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[11][24].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[11][25].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[11][25].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[11][25].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[11][25].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[11][25].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[11][25].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[11][25].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[11][25].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[11][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[11][25].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[11][26].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[11][26].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[11][26].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[11][26].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[11][26].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[11][26].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[11][26].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[11][26].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[11][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[11][26].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[11][27].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[11][27].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[11][27].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[11][27].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[11][27].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[11][27].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[11][27].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[11][27].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[11][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[11][27].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[11][28].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[11][28].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[11][28].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[11][28].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[11][28].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[11][28].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[11][28].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[11][28].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[11][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[11][28].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[11][29].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[11][29].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[11][29].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[11][29].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[11][29].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[11][29].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[11][29].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[11][29].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[11][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[11][29].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[11][30].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[11][30].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[11][30].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[11][30].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[11][30].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[11][30].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[11][30].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[11][30].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[11][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[11][30].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[11][31].dma__memc__write_valid      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[11][31].dma__memc__write_address    = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[11][31].dma__memc__write_data       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[11][31].dma__memc__read_valid       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[11][31].dma__memc__read_address     = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[11][31].dma__memc__read_pause       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[11][31].memc__dma__write_ready      = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[11][31].memc__dma__read_data        = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[11][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[11][31].memc__dma__read_ready       = pe_array_inst.pe_inst[11].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 12
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[12][0].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[12][0].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[12][0].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[12][0].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[12][0].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[12][0].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[12][0].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[12][0].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[12][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[12][0].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[12][1].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[12][1].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[12][1].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[12][1].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[12][1].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[12][1].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[12][1].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[12][1].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[12][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[12][1].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[12][2].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[12][2].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[12][2].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[12][2].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[12][2].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[12][2].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[12][2].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[12][2].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[12][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[12][2].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[12][3].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[12][3].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[12][3].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[12][3].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[12][3].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[12][3].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[12][3].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[12][3].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[12][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[12][3].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[12][4].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[12][4].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[12][4].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[12][4].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[12][4].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[12][4].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[12][4].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[12][4].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[12][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[12][4].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[12][5].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[12][5].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[12][5].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[12][5].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[12][5].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[12][5].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[12][5].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[12][5].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[12][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[12][5].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[12][6].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[12][6].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[12][6].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[12][6].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[12][6].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[12][6].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[12][6].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[12][6].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[12][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[12][6].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[12][7].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[12][7].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[12][7].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[12][7].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[12][7].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[12][7].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[12][7].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[12][7].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[12][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[12][7].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[12][8].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[12][8].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[12][8].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[12][8].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[12][8].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[12][8].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[12][8].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[12][8].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[12][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[12][8].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[12][9].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[12][9].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[12][9].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[12][9].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[12][9].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[12][9].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[12][9].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[12][9].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[12][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[12][9].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[12][10].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[12][10].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[12][10].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[12][10].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[12][10].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[12][10].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[12][10].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[12][10].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[12][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[12][10].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[12][11].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[12][11].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[12][11].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[12][11].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[12][11].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[12][11].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[12][11].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[12][11].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[12][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[12][11].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[12][12].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[12][12].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[12][12].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[12][12].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[12][12].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[12][12].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[12][12].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[12][12].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[12][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[12][12].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[12][13].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[12][13].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[12][13].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[12][13].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[12][13].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[12][13].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[12][13].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[12][13].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[12][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[12][13].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[12][14].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[12][14].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[12][14].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[12][14].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[12][14].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[12][14].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[12][14].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[12][14].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[12][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[12][14].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[12][15].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[12][15].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[12][15].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[12][15].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[12][15].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[12][15].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[12][15].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[12][15].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[12][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[12][15].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[12][16].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[12][16].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[12][16].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[12][16].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[12][16].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[12][16].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[12][16].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[12][16].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[12][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[12][16].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[12][17].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[12][17].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[12][17].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[12][17].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[12][17].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[12][17].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[12][17].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[12][17].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[12][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[12][17].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[12][18].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[12][18].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[12][18].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[12][18].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[12][18].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[12][18].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[12][18].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[12][18].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[12][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[12][18].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[12][19].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[12][19].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[12][19].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[12][19].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[12][19].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[12][19].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[12][19].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[12][19].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[12][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[12][19].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[12][20].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[12][20].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[12][20].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[12][20].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[12][20].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[12][20].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[12][20].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[12][20].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[12][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[12][20].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[12][21].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[12][21].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[12][21].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[12][21].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[12][21].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[12][21].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[12][21].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[12][21].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[12][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[12][21].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[12][22].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[12][22].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[12][22].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[12][22].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[12][22].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[12][22].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[12][22].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[12][22].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[12][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[12][22].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[12][23].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[12][23].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[12][23].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[12][23].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[12][23].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[12][23].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[12][23].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[12][23].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[12][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[12][23].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[12][24].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[12][24].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[12][24].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[12][24].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[12][24].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[12][24].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[12][24].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[12][24].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[12][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[12][24].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[12][25].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[12][25].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[12][25].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[12][25].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[12][25].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[12][25].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[12][25].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[12][25].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[12][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[12][25].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[12][26].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[12][26].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[12][26].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[12][26].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[12][26].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[12][26].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[12][26].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[12][26].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[12][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[12][26].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[12][27].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[12][27].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[12][27].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[12][27].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[12][27].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[12][27].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[12][27].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[12][27].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[12][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[12][27].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[12][28].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[12][28].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[12][28].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[12][28].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[12][28].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[12][28].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[12][28].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[12][28].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[12][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[12][28].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[12][29].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[12][29].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[12][29].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[12][29].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[12][29].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[12][29].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[12][29].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[12][29].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[12][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[12][29].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[12][30].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[12][30].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[12][30].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[12][30].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[12][30].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[12][30].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[12][30].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[12][30].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[12][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[12][30].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[12][31].dma__memc__write_valid      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[12][31].dma__memc__write_address    = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[12][31].dma__memc__write_data       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[12][31].dma__memc__read_valid       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[12][31].dma__memc__read_address     = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[12][31].dma__memc__read_pause       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[12][31].memc__dma__write_ready      = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[12][31].memc__dma__read_data        = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[12][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[12][31].memc__dma__read_ready       = pe_array_inst.pe_inst[12].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 13
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[13][0].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[13][0].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[13][0].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[13][0].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[13][0].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[13][0].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[13][0].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[13][0].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[13][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[13][0].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[13][1].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[13][1].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[13][1].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[13][1].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[13][1].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[13][1].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[13][1].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[13][1].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[13][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[13][1].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[13][2].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[13][2].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[13][2].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[13][2].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[13][2].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[13][2].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[13][2].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[13][2].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[13][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[13][2].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[13][3].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[13][3].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[13][3].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[13][3].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[13][3].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[13][3].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[13][3].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[13][3].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[13][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[13][3].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[13][4].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[13][4].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[13][4].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[13][4].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[13][4].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[13][4].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[13][4].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[13][4].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[13][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[13][4].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[13][5].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[13][5].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[13][5].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[13][5].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[13][5].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[13][5].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[13][5].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[13][5].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[13][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[13][5].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[13][6].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[13][6].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[13][6].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[13][6].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[13][6].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[13][6].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[13][6].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[13][6].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[13][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[13][6].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[13][7].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[13][7].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[13][7].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[13][7].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[13][7].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[13][7].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[13][7].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[13][7].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[13][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[13][7].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[13][8].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[13][8].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[13][8].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[13][8].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[13][8].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[13][8].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[13][8].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[13][8].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[13][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[13][8].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[13][9].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[13][9].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[13][9].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[13][9].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[13][9].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[13][9].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[13][9].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[13][9].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[13][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[13][9].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[13][10].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[13][10].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[13][10].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[13][10].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[13][10].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[13][10].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[13][10].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[13][10].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[13][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[13][10].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[13][11].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[13][11].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[13][11].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[13][11].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[13][11].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[13][11].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[13][11].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[13][11].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[13][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[13][11].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[13][12].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[13][12].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[13][12].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[13][12].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[13][12].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[13][12].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[13][12].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[13][12].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[13][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[13][12].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[13][13].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[13][13].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[13][13].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[13][13].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[13][13].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[13][13].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[13][13].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[13][13].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[13][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[13][13].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[13][14].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[13][14].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[13][14].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[13][14].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[13][14].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[13][14].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[13][14].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[13][14].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[13][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[13][14].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[13][15].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[13][15].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[13][15].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[13][15].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[13][15].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[13][15].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[13][15].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[13][15].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[13][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[13][15].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[13][16].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[13][16].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[13][16].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[13][16].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[13][16].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[13][16].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[13][16].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[13][16].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[13][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[13][16].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[13][17].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[13][17].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[13][17].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[13][17].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[13][17].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[13][17].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[13][17].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[13][17].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[13][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[13][17].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[13][18].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[13][18].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[13][18].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[13][18].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[13][18].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[13][18].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[13][18].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[13][18].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[13][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[13][18].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[13][19].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[13][19].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[13][19].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[13][19].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[13][19].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[13][19].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[13][19].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[13][19].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[13][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[13][19].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[13][20].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[13][20].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[13][20].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[13][20].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[13][20].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[13][20].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[13][20].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[13][20].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[13][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[13][20].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[13][21].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[13][21].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[13][21].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[13][21].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[13][21].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[13][21].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[13][21].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[13][21].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[13][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[13][21].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[13][22].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[13][22].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[13][22].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[13][22].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[13][22].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[13][22].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[13][22].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[13][22].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[13][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[13][22].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[13][23].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[13][23].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[13][23].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[13][23].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[13][23].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[13][23].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[13][23].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[13][23].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[13][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[13][23].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[13][24].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[13][24].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[13][24].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[13][24].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[13][24].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[13][24].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[13][24].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[13][24].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[13][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[13][24].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[13][25].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[13][25].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[13][25].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[13][25].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[13][25].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[13][25].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[13][25].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[13][25].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[13][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[13][25].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[13][26].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[13][26].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[13][26].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[13][26].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[13][26].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[13][26].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[13][26].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[13][26].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[13][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[13][26].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[13][27].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[13][27].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[13][27].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[13][27].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[13][27].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[13][27].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[13][27].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[13][27].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[13][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[13][27].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[13][28].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[13][28].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[13][28].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[13][28].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[13][28].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[13][28].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[13][28].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[13][28].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[13][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[13][28].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[13][29].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[13][29].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[13][29].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[13][29].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[13][29].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[13][29].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[13][29].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[13][29].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[13][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[13][29].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[13][30].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[13][30].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[13][30].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[13][30].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[13][30].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[13][30].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[13][30].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[13][30].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[13][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[13][30].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[13][31].dma__memc__write_valid      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[13][31].dma__memc__write_address    = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[13][31].dma__memc__write_data       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[13][31].dma__memc__read_valid       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[13][31].dma__memc__read_address     = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[13][31].dma__memc__read_pause       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[13][31].memc__dma__write_ready      = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[13][31].memc__dma__read_data        = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[13][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[13][31].memc__dma__read_ready       = pe_array_inst.pe_inst[13].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 14
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[14][0].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[14][0].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[14][0].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[14][0].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[14][0].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[14][0].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[14][0].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[14][0].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[14][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[14][0].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[14][1].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[14][1].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[14][1].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[14][1].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[14][1].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[14][1].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[14][1].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[14][1].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[14][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[14][1].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[14][2].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[14][2].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[14][2].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[14][2].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[14][2].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[14][2].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[14][2].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[14][2].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[14][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[14][2].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[14][3].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[14][3].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[14][3].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[14][3].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[14][3].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[14][3].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[14][3].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[14][3].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[14][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[14][3].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[14][4].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[14][4].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[14][4].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[14][4].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[14][4].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[14][4].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[14][4].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[14][4].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[14][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[14][4].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[14][5].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[14][5].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[14][5].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[14][5].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[14][5].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[14][5].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[14][5].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[14][5].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[14][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[14][5].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[14][6].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[14][6].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[14][6].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[14][6].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[14][6].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[14][6].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[14][6].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[14][6].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[14][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[14][6].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[14][7].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[14][7].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[14][7].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[14][7].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[14][7].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[14][7].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[14][7].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[14][7].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[14][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[14][7].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[14][8].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[14][8].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[14][8].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[14][8].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[14][8].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[14][8].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[14][8].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[14][8].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[14][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[14][8].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[14][9].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[14][9].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[14][9].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[14][9].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[14][9].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[14][9].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[14][9].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[14][9].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[14][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[14][9].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[14][10].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[14][10].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[14][10].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[14][10].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[14][10].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[14][10].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[14][10].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[14][10].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[14][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[14][10].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[14][11].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[14][11].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[14][11].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[14][11].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[14][11].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[14][11].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[14][11].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[14][11].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[14][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[14][11].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[14][12].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[14][12].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[14][12].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[14][12].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[14][12].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[14][12].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[14][12].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[14][12].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[14][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[14][12].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[14][13].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[14][13].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[14][13].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[14][13].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[14][13].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[14][13].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[14][13].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[14][13].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[14][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[14][13].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[14][14].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[14][14].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[14][14].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[14][14].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[14][14].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[14][14].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[14][14].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[14][14].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[14][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[14][14].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[14][15].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[14][15].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[14][15].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[14][15].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[14][15].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[14][15].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[14][15].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[14][15].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[14][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[14][15].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[14][16].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[14][16].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[14][16].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[14][16].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[14][16].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[14][16].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[14][16].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[14][16].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[14][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[14][16].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[14][17].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[14][17].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[14][17].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[14][17].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[14][17].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[14][17].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[14][17].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[14][17].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[14][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[14][17].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[14][18].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[14][18].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[14][18].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[14][18].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[14][18].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[14][18].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[14][18].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[14][18].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[14][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[14][18].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[14][19].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[14][19].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[14][19].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[14][19].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[14][19].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[14][19].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[14][19].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[14][19].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[14][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[14][19].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[14][20].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[14][20].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[14][20].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[14][20].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[14][20].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[14][20].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[14][20].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[14][20].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[14][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[14][20].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[14][21].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[14][21].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[14][21].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[14][21].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[14][21].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[14][21].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[14][21].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[14][21].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[14][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[14][21].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[14][22].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[14][22].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[14][22].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[14][22].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[14][22].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[14][22].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[14][22].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[14][22].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[14][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[14][22].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[14][23].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[14][23].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[14][23].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[14][23].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[14][23].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[14][23].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[14][23].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[14][23].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[14][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[14][23].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[14][24].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[14][24].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[14][24].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[14][24].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[14][24].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[14][24].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[14][24].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[14][24].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[14][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[14][24].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[14][25].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[14][25].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[14][25].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[14][25].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[14][25].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[14][25].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[14][25].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[14][25].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[14][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[14][25].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[14][26].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[14][26].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[14][26].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[14][26].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[14][26].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[14][26].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[14][26].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[14][26].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[14][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[14][26].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[14][27].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[14][27].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[14][27].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[14][27].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[14][27].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[14][27].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[14][27].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[14][27].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[14][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[14][27].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[14][28].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[14][28].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[14][28].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[14][28].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[14][28].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[14][28].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[14][28].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[14][28].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[14][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[14][28].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[14][29].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[14][29].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[14][29].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[14][29].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[14][29].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[14][29].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[14][29].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[14][29].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[14][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[14][29].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[14][30].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[14][30].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[14][30].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[14][30].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[14][30].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[14][30].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[14][30].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[14][30].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[14][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[14][30].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[14][31].dma__memc__write_valid      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[14][31].dma__memc__write_address    = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[14][31].dma__memc__write_data       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[14][31].dma__memc__read_valid       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[14][31].dma__memc__read_address     = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[14][31].dma__memc__read_pause       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[14][31].memc__dma__write_ready      = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[14][31].memc__dma__read_data        = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[14][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[14][31].memc__dma__read_ready       = pe_array_inst.pe_inst[14].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 15
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[15][0].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[15][0].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[15][0].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[15][0].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[15][0].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[15][0].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[15][0].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[15][0].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[15][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[15][0].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[15][1].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[15][1].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[15][1].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[15][1].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[15][1].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[15][1].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[15][1].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[15][1].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[15][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[15][1].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[15][2].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[15][2].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[15][2].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[15][2].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[15][2].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[15][2].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[15][2].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[15][2].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[15][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[15][2].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[15][3].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[15][3].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[15][3].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[15][3].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[15][3].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[15][3].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[15][3].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[15][3].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[15][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[15][3].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[15][4].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[15][4].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[15][4].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[15][4].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[15][4].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[15][4].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[15][4].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[15][4].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[15][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[15][4].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[15][5].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[15][5].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[15][5].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[15][5].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[15][5].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[15][5].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[15][5].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[15][5].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[15][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[15][5].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[15][6].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[15][6].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[15][6].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[15][6].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[15][6].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[15][6].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[15][6].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[15][6].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[15][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[15][6].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[15][7].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[15][7].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[15][7].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[15][7].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[15][7].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[15][7].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[15][7].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[15][7].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[15][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[15][7].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[15][8].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[15][8].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[15][8].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[15][8].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[15][8].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[15][8].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[15][8].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[15][8].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[15][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[15][8].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[15][9].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[15][9].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[15][9].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[15][9].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[15][9].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[15][9].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[15][9].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[15][9].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[15][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[15][9].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[15][10].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[15][10].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[15][10].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[15][10].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[15][10].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[15][10].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[15][10].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[15][10].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[15][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[15][10].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[15][11].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[15][11].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[15][11].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[15][11].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[15][11].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[15][11].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[15][11].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[15][11].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[15][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[15][11].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[15][12].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[15][12].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[15][12].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[15][12].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[15][12].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[15][12].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[15][12].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[15][12].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[15][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[15][12].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[15][13].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[15][13].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[15][13].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[15][13].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[15][13].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[15][13].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[15][13].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[15][13].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[15][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[15][13].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[15][14].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[15][14].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[15][14].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[15][14].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[15][14].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[15][14].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[15][14].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[15][14].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[15][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[15][14].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[15][15].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[15][15].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[15][15].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[15][15].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[15][15].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[15][15].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[15][15].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[15][15].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[15][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[15][15].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[15][16].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[15][16].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[15][16].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[15][16].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[15][16].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[15][16].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[15][16].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[15][16].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[15][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[15][16].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[15][17].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[15][17].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[15][17].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[15][17].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[15][17].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[15][17].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[15][17].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[15][17].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[15][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[15][17].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[15][18].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[15][18].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[15][18].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[15][18].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[15][18].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[15][18].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[15][18].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[15][18].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[15][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[15][18].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[15][19].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[15][19].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[15][19].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[15][19].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[15][19].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[15][19].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[15][19].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[15][19].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[15][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[15][19].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[15][20].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[15][20].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[15][20].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[15][20].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[15][20].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[15][20].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[15][20].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[15][20].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[15][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[15][20].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[15][21].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[15][21].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[15][21].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[15][21].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[15][21].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[15][21].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[15][21].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[15][21].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[15][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[15][21].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[15][22].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[15][22].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[15][22].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[15][22].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[15][22].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[15][22].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[15][22].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[15][22].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[15][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[15][22].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[15][23].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[15][23].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[15][23].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[15][23].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[15][23].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[15][23].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[15][23].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[15][23].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[15][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[15][23].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[15][24].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[15][24].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[15][24].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[15][24].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[15][24].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[15][24].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[15][24].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[15][24].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[15][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[15][24].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[15][25].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[15][25].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[15][25].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[15][25].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[15][25].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[15][25].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[15][25].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[15][25].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[15][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[15][25].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[15][26].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[15][26].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[15][26].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[15][26].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[15][26].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[15][26].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[15][26].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[15][26].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[15][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[15][26].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[15][27].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[15][27].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[15][27].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[15][27].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[15][27].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[15][27].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[15][27].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[15][27].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[15][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[15][27].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[15][28].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[15][28].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[15][28].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[15][28].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[15][28].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[15][28].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[15][28].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[15][28].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[15][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[15][28].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[15][29].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[15][29].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[15][29].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[15][29].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[15][29].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[15][29].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[15][29].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[15][29].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[15][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[15][29].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[15][30].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[15][30].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[15][30].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[15][30].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[15][30].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[15][30].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[15][30].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[15][30].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[15][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[15][30].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[15][31].dma__memc__write_valid      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[15][31].dma__memc__write_address    = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[15][31].dma__memc__write_data       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[15][31].dma__memc__read_valid       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[15][31].dma__memc__read_address     = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[15][31].dma__memc__read_pause       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[15][31].memc__dma__write_ready      = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[15][31].memc__dma__read_data        = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[15][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[15][31].memc__dma__read_ready       = pe_array_inst.pe_inst[15].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 16
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[16][0].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[16][0].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[16][0].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[16][0].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[16][0].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[16][0].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[16][0].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[16][0].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[16][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[16][0].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[16][1].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[16][1].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[16][1].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[16][1].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[16][1].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[16][1].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[16][1].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[16][1].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[16][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[16][1].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[16][2].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[16][2].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[16][2].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[16][2].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[16][2].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[16][2].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[16][2].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[16][2].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[16][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[16][2].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[16][3].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[16][3].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[16][3].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[16][3].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[16][3].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[16][3].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[16][3].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[16][3].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[16][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[16][3].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[16][4].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[16][4].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[16][4].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[16][4].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[16][4].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[16][4].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[16][4].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[16][4].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[16][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[16][4].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[16][5].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[16][5].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[16][5].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[16][5].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[16][5].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[16][5].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[16][5].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[16][5].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[16][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[16][5].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[16][6].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[16][6].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[16][6].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[16][6].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[16][6].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[16][6].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[16][6].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[16][6].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[16][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[16][6].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[16][7].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[16][7].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[16][7].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[16][7].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[16][7].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[16][7].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[16][7].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[16][7].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[16][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[16][7].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[16][8].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[16][8].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[16][8].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[16][8].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[16][8].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[16][8].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[16][8].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[16][8].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[16][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[16][8].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[16][9].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[16][9].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[16][9].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[16][9].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[16][9].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[16][9].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[16][9].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[16][9].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[16][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[16][9].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[16][10].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[16][10].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[16][10].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[16][10].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[16][10].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[16][10].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[16][10].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[16][10].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[16][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[16][10].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[16][11].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[16][11].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[16][11].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[16][11].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[16][11].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[16][11].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[16][11].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[16][11].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[16][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[16][11].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[16][12].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[16][12].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[16][12].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[16][12].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[16][12].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[16][12].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[16][12].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[16][12].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[16][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[16][12].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[16][13].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[16][13].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[16][13].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[16][13].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[16][13].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[16][13].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[16][13].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[16][13].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[16][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[16][13].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[16][14].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[16][14].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[16][14].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[16][14].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[16][14].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[16][14].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[16][14].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[16][14].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[16][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[16][14].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[16][15].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[16][15].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[16][15].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[16][15].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[16][15].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[16][15].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[16][15].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[16][15].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[16][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[16][15].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[16][16].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[16][16].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[16][16].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[16][16].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[16][16].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[16][16].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[16][16].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[16][16].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[16][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[16][16].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[16][17].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[16][17].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[16][17].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[16][17].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[16][17].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[16][17].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[16][17].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[16][17].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[16][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[16][17].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[16][18].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[16][18].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[16][18].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[16][18].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[16][18].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[16][18].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[16][18].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[16][18].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[16][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[16][18].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[16][19].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[16][19].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[16][19].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[16][19].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[16][19].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[16][19].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[16][19].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[16][19].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[16][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[16][19].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[16][20].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[16][20].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[16][20].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[16][20].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[16][20].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[16][20].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[16][20].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[16][20].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[16][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[16][20].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[16][21].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[16][21].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[16][21].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[16][21].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[16][21].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[16][21].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[16][21].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[16][21].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[16][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[16][21].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[16][22].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[16][22].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[16][22].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[16][22].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[16][22].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[16][22].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[16][22].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[16][22].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[16][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[16][22].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[16][23].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[16][23].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[16][23].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[16][23].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[16][23].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[16][23].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[16][23].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[16][23].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[16][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[16][23].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[16][24].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[16][24].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[16][24].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[16][24].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[16][24].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[16][24].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[16][24].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[16][24].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[16][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[16][24].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[16][25].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[16][25].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[16][25].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[16][25].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[16][25].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[16][25].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[16][25].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[16][25].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[16][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[16][25].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[16][26].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[16][26].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[16][26].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[16][26].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[16][26].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[16][26].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[16][26].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[16][26].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[16][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[16][26].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[16][27].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[16][27].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[16][27].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[16][27].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[16][27].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[16][27].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[16][27].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[16][27].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[16][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[16][27].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[16][28].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[16][28].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[16][28].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[16][28].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[16][28].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[16][28].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[16][28].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[16][28].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[16][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[16][28].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[16][29].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[16][29].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[16][29].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[16][29].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[16][29].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[16][29].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[16][29].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[16][29].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[16][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[16][29].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[16][30].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[16][30].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[16][30].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[16][30].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[16][30].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[16][30].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[16][30].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[16][30].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[16][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[16][30].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[16][31].dma__memc__write_valid      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[16][31].dma__memc__write_address    = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[16][31].dma__memc__write_data       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[16][31].dma__memc__read_valid       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[16][31].dma__memc__read_address     = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[16][31].dma__memc__read_pause       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[16][31].memc__dma__write_ready      = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[16][31].memc__dma__read_data        = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[16][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[16][31].memc__dma__read_ready       = pe_array_inst.pe_inst[16].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 17
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[17][0].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[17][0].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[17][0].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[17][0].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[17][0].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[17][0].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[17][0].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[17][0].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[17][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[17][0].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[17][1].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[17][1].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[17][1].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[17][1].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[17][1].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[17][1].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[17][1].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[17][1].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[17][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[17][1].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[17][2].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[17][2].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[17][2].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[17][2].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[17][2].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[17][2].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[17][2].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[17][2].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[17][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[17][2].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[17][3].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[17][3].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[17][3].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[17][3].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[17][3].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[17][3].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[17][3].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[17][3].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[17][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[17][3].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[17][4].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[17][4].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[17][4].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[17][4].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[17][4].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[17][4].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[17][4].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[17][4].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[17][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[17][4].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[17][5].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[17][5].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[17][5].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[17][5].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[17][5].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[17][5].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[17][5].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[17][5].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[17][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[17][5].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[17][6].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[17][6].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[17][6].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[17][6].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[17][6].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[17][6].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[17][6].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[17][6].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[17][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[17][6].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[17][7].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[17][7].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[17][7].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[17][7].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[17][7].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[17][7].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[17][7].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[17][7].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[17][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[17][7].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[17][8].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[17][8].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[17][8].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[17][8].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[17][8].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[17][8].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[17][8].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[17][8].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[17][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[17][8].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[17][9].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[17][9].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[17][9].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[17][9].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[17][9].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[17][9].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[17][9].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[17][9].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[17][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[17][9].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[17][10].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[17][10].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[17][10].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[17][10].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[17][10].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[17][10].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[17][10].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[17][10].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[17][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[17][10].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[17][11].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[17][11].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[17][11].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[17][11].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[17][11].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[17][11].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[17][11].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[17][11].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[17][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[17][11].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[17][12].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[17][12].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[17][12].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[17][12].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[17][12].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[17][12].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[17][12].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[17][12].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[17][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[17][12].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[17][13].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[17][13].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[17][13].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[17][13].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[17][13].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[17][13].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[17][13].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[17][13].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[17][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[17][13].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[17][14].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[17][14].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[17][14].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[17][14].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[17][14].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[17][14].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[17][14].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[17][14].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[17][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[17][14].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[17][15].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[17][15].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[17][15].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[17][15].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[17][15].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[17][15].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[17][15].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[17][15].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[17][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[17][15].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[17][16].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[17][16].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[17][16].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[17][16].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[17][16].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[17][16].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[17][16].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[17][16].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[17][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[17][16].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[17][17].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[17][17].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[17][17].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[17][17].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[17][17].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[17][17].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[17][17].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[17][17].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[17][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[17][17].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[17][18].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[17][18].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[17][18].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[17][18].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[17][18].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[17][18].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[17][18].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[17][18].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[17][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[17][18].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[17][19].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[17][19].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[17][19].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[17][19].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[17][19].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[17][19].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[17][19].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[17][19].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[17][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[17][19].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[17][20].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[17][20].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[17][20].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[17][20].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[17][20].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[17][20].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[17][20].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[17][20].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[17][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[17][20].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[17][21].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[17][21].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[17][21].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[17][21].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[17][21].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[17][21].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[17][21].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[17][21].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[17][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[17][21].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[17][22].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[17][22].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[17][22].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[17][22].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[17][22].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[17][22].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[17][22].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[17][22].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[17][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[17][22].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[17][23].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[17][23].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[17][23].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[17][23].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[17][23].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[17][23].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[17][23].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[17][23].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[17][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[17][23].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[17][24].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[17][24].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[17][24].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[17][24].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[17][24].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[17][24].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[17][24].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[17][24].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[17][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[17][24].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[17][25].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[17][25].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[17][25].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[17][25].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[17][25].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[17][25].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[17][25].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[17][25].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[17][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[17][25].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[17][26].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[17][26].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[17][26].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[17][26].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[17][26].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[17][26].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[17][26].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[17][26].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[17][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[17][26].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[17][27].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[17][27].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[17][27].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[17][27].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[17][27].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[17][27].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[17][27].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[17][27].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[17][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[17][27].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[17][28].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[17][28].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[17][28].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[17][28].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[17][28].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[17][28].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[17][28].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[17][28].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[17][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[17][28].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[17][29].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[17][29].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[17][29].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[17][29].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[17][29].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[17][29].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[17][29].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[17][29].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[17][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[17][29].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[17][30].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[17][30].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[17][30].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[17][30].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[17][30].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[17][30].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[17][30].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[17][30].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[17][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[17][30].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[17][31].dma__memc__write_valid      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[17][31].dma__memc__write_address    = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[17][31].dma__memc__write_data       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[17][31].dma__memc__read_valid       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[17][31].dma__memc__read_address     = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[17][31].dma__memc__read_pause       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[17][31].memc__dma__write_ready      = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[17][31].memc__dma__read_data        = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[17][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[17][31].memc__dma__read_ready       = pe_array_inst.pe_inst[17].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 18
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[18][0].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[18][0].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[18][0].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[18][0].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[18][0].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[18][0].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[18][0].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[18][0].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[18][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[18][0].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[18][1].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[18][1].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[18][1].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[18][1].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[18][1].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[18][1].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[18][1].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[18][1].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[18][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[18][1].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[18][2].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[18][2].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[18][2].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[18][2].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[18][2].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[18][2].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[18][2].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[18][2].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[18][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[18][2].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[18][3].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[18][3].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[18][3].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[18][3].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[18][3].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[18][3].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[18][3].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[18][3].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[18][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[18][3].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[18][4].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[18][4].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[18][4].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[18][4].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[18][4].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[18][4].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[18][4].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[18][4].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[18][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[18][4].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[18][5].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[18][5].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[18][5].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[18][5].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[18][5].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[18][5].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[18][5].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[18][5].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[18][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[18][5].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[18][6].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[18][6].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[18][6].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[18][6].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[18][6].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[18][6].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[18][6].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[18][6].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[18][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[18][6].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[18][7].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[18][7].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[18][7].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[18][7].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[18][7].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[18][7].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[18][7].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[18][7].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[18][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[18][7].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[18][8].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[18][8].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[18][8].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[18][8].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[18][8].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[18][8].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[18][8].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[18][8].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[18][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[18][8].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[18][9].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[18][9].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[18][9].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[18][9].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[18][9].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[18][9].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[18][9].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[18][9].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[18][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[18][9].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[18][10].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[18][10].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[18][10].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[18][10].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[18][10].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[18][10].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[18][10].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[18][10].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[18][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[18][10].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[18][11].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[18][11].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[18][11].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[18][11].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[18][11].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[18][11].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[18][11].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[18][11].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[18][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[18][11].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[18][12].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[18][12].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[18][12].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[18][12].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[18][12].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[18][12].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[18][12].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[18][12].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[18][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[18][12].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[18][13].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[18][13].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[18][13].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[18][13].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[18][13].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[18][13].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[18][13].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[18][13].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[18][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[18][13].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[18][14].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[18][14].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[18][14].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[18][14].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[18][14].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[18][14].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[18][14].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[18][14].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[18][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[18][14].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[18][15].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[18][15].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[18][15].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[18][15].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[18][15].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[18][15].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[18][15].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[18][15].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[18][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[18][15].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[18][16].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[18][16].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[18][16].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[18][16].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[18][16].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[18][16].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[18][16].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[18][16].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[18][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[18][16].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[18][17].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[18][17].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[18][17].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[18][17].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[18][17].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[18][17].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[18][17].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[18][17].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[18][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[18][17].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[18][18].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[18][18].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[18][18].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[18][18].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[18][18].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[18][18].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[18][18].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[18][18].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[18][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[18][18].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[18][19].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[18][19].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[18][19].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[18][19].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[18][19].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[18][19].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[18][19].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[18][19].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[18][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[18][19].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[18][20].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[18][20].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[18][20].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[18][20].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[18][20].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[18][20].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[18][20].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[18][20].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[18][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[18][20].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[18][21].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[18][21].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[18][21].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[18][21].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[18][21].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[18][21].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[18][21].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[18][21].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[18][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[18][21].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[18][22].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[18][22].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[18][22].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[18][22].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[18][22].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[18][22].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[18][22].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[18][22].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[18][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[18][22].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[18][23].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[18][23].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[18][23].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[18][23].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[18][23].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[18][23].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[18][23].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[18][23].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[18][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[18][23].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[18][24].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[18][24].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[18][24].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[18][24].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[18][24].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[18][24].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[18][24].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[18][24].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[18][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[18][24].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[18][25].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[18][25].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[18][25].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[18][25].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[18][25].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[18][25].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[18][25].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[18][25].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[18][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[18][25].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[18][26].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[18][26].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[18][26].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[18][26].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[18][26].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[18][26].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[18][26].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[18][26].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[18][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[18][26].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[18][27].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[18][27].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[18][27].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[18][27].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[18][27].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[18][27].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[18][27].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[18][27].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[18][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[18][27].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[18][28].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[18][28].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[18][28].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[18][28].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[18][28].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[18][28].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[18][28].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[18][28].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[18][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[18][28].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[18][29].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[18][29].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[18][29].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[18][29].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[18][29].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[18][29].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[18][29].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[18][29].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[18][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[18][29].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[18][30].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[18][30].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[18][30].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[18][30].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[18][30].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[18][30].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[18][30].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[18][30].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[18][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[18][30].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[18][31].dma__memc__write_valid      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[18][31].dma__memc__write_address    = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[18][31].dma__memc__write_data       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[18][31].dma__memc__read_valid       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[18][31].dma__memc__read_address     = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[18][31].dma__memc__read_pause       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[18][31].memc__dma__write_ready      = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[18][31].memc__dma__read_data        = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[18][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[18][31].memc__dma__read_ready       = pe_array_inst.pe_inst[18].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 19
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[19][0].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[19][0].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[19][0].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[19][0].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[19][0].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[19][0].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[19][0].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[19][0].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[19][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[19][0].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[19][1].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[19][1].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[19][1].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[19][1].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[19][1].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[19][1].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[19][1].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[19][1].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[19][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[19][1].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[19][2].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[19][2].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[19][2].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[19][2].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[19][2].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[19][2].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[19][2].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[19][2].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[19][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[19][2].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[19][3].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[19][3].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[19][3].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[19][3].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[19][3].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[19][3].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[19][3].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[19][3].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[19][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[19][3].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[19][4].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[19][4].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[19][4].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[19][4].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[19][4].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[19][4].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[19][4].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[19][4].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[19][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[19][4].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[19][5].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[19][5].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[19][5].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[19][5].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[19][5].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[19][5].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[19][5].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[19][5].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[19][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[19][5].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[19][6].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[19][6].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[19][6].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[19][6].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[19][6].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[19][6].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[19][6].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[19][6].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[19][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[19][6].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[19][7].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[19][7].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[19][7].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[19][7].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[19][7].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[19][7].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[19][7].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[19][7].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[19][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[19][7].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[19][8].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[19][8].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[19][8].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[19][8].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[19][8].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[19][8].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[19][8].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[19][8].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[19][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[19][8].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[19][9].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[19][9].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[19][9].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[19][9].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[19][9].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[19][9].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[19][9].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[19][9].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[19][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[19][9].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[19][10].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[19][10].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[19][10].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[19][10].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[19][10].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[19][10].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[19][10].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[19][10].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[19][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[19][10].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[19][11].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[19][11].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[19][11].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[19][11].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[19][11].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[19][11].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[19][11].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[19][11].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[19][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[19][11].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[19][12].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[19][12].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[19][12].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[19][12].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[19][12].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[19][12].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[19][12].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[19][12].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[19][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[19][12].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[19][13].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[19][13].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[19][13].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[19][13].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[19][13].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[19][13].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[19][13].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[19][13].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[19][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[19][13].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[19][14].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[19][14].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[19][14].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[19][14].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[19][14].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[19][14].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[19][14].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[19][14].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[19][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[19][14].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[19][15].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[19][15].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[19][15].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[19][15].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[19][15].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[19][15].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[19][15].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[19][15].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[19][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[19][15].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[19][16].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[19][16].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[19][16].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[19][16].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[19][16].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[19][16].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[19][16].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[19][16].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[19][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[19][16].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[19][17].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[19][17].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[19][17].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[19][17].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[19][17].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[19][17].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[19][17].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[19][17].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[19][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[19][17].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[19][18].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[19][18].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[19][18].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[19][18].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[19][18].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[19][18].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[19][18].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[19][18].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[19][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[19][18].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[19][19].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[19][19].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[19][19].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[19][19].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[19][19].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[19][19].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[19][19].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[19][19].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[19][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[19][19].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[19][20].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[19][20].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[19][20].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[19][20].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[19][20].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[19][20].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[19][20].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[19][20].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[19][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[19][20].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[19][21].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[19][21].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[19][21].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[19][21].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[19][21].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[19][21].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[19][21].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[19][21].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[19][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[19][21].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[19][22].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[19][22].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[19][22].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[19][22].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[19][22].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[19][22].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[19][22].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[19][22].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[19][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[19][22].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[19][23].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[19][23].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[19][23].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[19][23].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[19][23].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[19][23].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[19][23].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[19][23].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[19][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[19][23].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[19][24].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[19][24].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[19][24].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[19][24].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[19][24].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[19][24].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[19][24].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[19][24].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[19][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[19][24].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[19][25].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[19][25].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[19][25].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[19][25].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[19][25].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[19][25].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[19][25].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[19][25].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[19][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[19][25].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[19][26].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[19][26].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[19][26].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[19][26].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[19][26].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[19][26].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[19][26].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[19][26].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[19][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[19][26].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[19][27].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[19][27].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[19][27].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[19][27].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[19][27].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[19][27].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[19][27].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[19][27].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[19][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[19][27].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[19][28].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[19][28].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[19][28].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[19][28].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[19][28].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[19][28].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[19][28].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[19][28].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[19][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[19][28].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[19][29].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[19][29].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[19][29].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[19][29].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[19][29].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[19][29].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[19][29].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[19][29].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[19][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[19][29].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[19][30].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[19][30].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[19][30].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[19][30].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[19][30].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[19][30].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[19][30].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[19][30].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[19][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[19][30].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[19][31].dma__memc__write_valid      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[19][31].dma__memc__write_address    = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[19][31].dma__memc__write_data       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[19][31].dma__memc__read_valid       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[19][31].dma__memc__read_address     = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[19][31].dma__memc__read_pause       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[19][31].memc__dma__write_ready      = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[19][31].memc__dma__read_data        = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[19][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[19][31].memc__dma__read_ready       = pe_array_inst.pe_inst[19].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 20
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[20][0].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[20][0].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[20][0].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[20][0].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[20][0].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[20][0].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[20][0].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[20][0].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[20][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[20][0].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[20][1].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[20][1].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[20][1].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[20][1].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[20][1].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[20][1].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[20][1].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[20][1].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[20][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[20][1].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[20][2].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[20][2].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[20][2].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[20][2].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[20][2].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[20][2].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[20][2].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[20][2].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[20][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[20][2].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[20][3].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[20][3].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[20][3].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[20][3].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[20][3].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[20][3].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[20][3].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[20][3].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[20][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[20][3].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[20][4].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[20][4].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[20][4].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[20][4].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[20][4].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[20][4].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[20][4].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[20][4].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[20][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[20][4].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[20][5].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[20][5].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[20][5].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[20][5].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[20][5].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[20][5].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[20][5].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[20][5].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[20][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[20][5].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[20][6].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[20][6].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[20][6].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[20][6].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[20][6].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[20][6].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[20][6].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[20][6].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[20][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[20][6].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[20][7].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[20][7].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[20][7].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[20][7].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[20][7].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[20][7].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[20][7].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[20][7].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[20][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[20][7].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[20][8].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[20][8].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[20][8].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[20][8].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[20][8].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[20][8].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[20][8].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[20][8].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[20][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[20][8].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[20][9].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[20][9].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[20][9].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[20][9].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[20][9].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[20][9].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[20][9].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[20][9].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[20][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[20][9].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[20][10].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[20][10].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[20][10].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[20][10].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[20][10].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[20][10].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[20][10].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[20][10].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[20][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[20][10].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[20][11].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[20][11].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[20][11].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[20][11].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[20][11].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[20][11].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[20][11].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[20][11].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[20][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[20][11].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[20][12].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[20][12].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[20][12].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[20][12].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[20][12].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[20][12].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[20][12].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[20][12].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[20][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[20][12].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[20][13].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[20][13].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[20][13].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[20][13].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[20][13].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[20][13].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[20][13].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[20][13].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[20][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[20][13].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[20][14].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[20][14].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[20][14].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[20][14].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[20][14].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[20][14].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[20][14].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[20][14].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[20][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[20][14].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[20][15].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[20][15].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[20][15].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[20][15].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[20][15].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[20][15].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[20][15].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[20][15].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[20][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[20][15].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[20][16].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[20][16].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[20][16].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[20][16].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[20][16].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[20][16].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[20][16].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[20][16].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[20][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[20][16].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[20][17].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[20][17].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[20][17].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[20][17].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[20][17].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[20][17].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[20][17].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[20][17].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[20][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[20][17].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[20][18].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[20][18].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[20][18].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[20][18].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[20][18].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[20][18].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[20][18].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[20][18].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[20][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[20][18].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[20][19].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[20][19].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[20][19].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[20][19].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[20][19].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[20][19].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[20][19].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[20][19].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[20][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[20][19].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[20][20].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[20][20].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[20][20].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[20][20].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[20][20].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[20][20].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[20][20].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[20][20].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[20][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[20][20].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[20][21].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[20][21].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[20][21].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[20][21].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[20][21].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[20][21].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[20][21].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[20][21].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[20][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[20][21].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[20][22].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[20][22].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[20][22].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[20][22].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[20][22].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[20][22].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[20][22].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[20][22].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[20][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[20][22].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[20][23].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[20][23].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[20][23].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[20][23].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[20][23].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[20][23].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[20][23].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[20][23].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[20][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[20][23].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[20][24].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[20][24].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[20][24].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[20][24].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[20][24].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[20][24].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[20][24].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[20][24].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[20][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[20][24].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[20][25].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[20][25].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[20][25].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[20][25].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[20][25].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[20][25].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[20][25].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[20][25].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[20][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[20][25].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[20][26].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[20][26].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[20][26].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[20][26].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[20][26].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[20][26].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[20][26].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[20][26].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[20][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[20][26].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[20][27].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[20][27].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[20][27].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[20][27].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[20][27].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[20][27].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[20][27].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[20][27].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[20][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[20][27].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[20][28].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[20][28].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[20][28].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[20][28].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[20][28].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[20][28].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[20][28].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[20][28].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[20][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[20][28].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[20][29].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[20][29].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[20][29].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[20][29].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[20][29].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[20][29].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[20][29].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[20][29].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[20][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[20][29].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[20][30].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[20][30].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[20][30].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[20][30].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[20][30].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[20][30].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[20][30].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[20][30].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[20][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[20][30].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[20][31].dma__memc__write_valid      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[20][31].dma__memc__write_address    = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[20][31].dma__memc__write_data       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[20][31].dma__memc__read_valid       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[20][31].dma__memc__read_address     = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[20][31].dma__memc__read_pause       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[20][31].memc__dma__write_ready      = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[20][31].memc__dma__read_data        = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[20][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[20][31].memc__dma__read_ready       = pe_array_inst.pe_inst[20].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 21
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[21][0].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[21][0].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[21][0].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[21][0].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[21][0].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[21][0].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[21][0].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[21][0].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[21][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[21][0].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[21][1].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[21][1].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[21][1].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[21][1].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[21][1].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[21][1].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[21][1].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[21][1].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[21][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[21][1].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[21][2].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[21][2].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[21][2].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[21][2].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[21][2].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[21][2].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[21][2].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[21][2].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[21][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[21][2].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[21][3].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[21][3].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[21][3].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[21][3].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[21][3].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[21][3].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[21][3].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[21][3].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[21][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[21][3].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[21][4].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[21][4].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[21][4].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[21][4].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[21][4].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[21][4].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[21][4].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[21][4].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[21][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[21][4].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[21][5].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[21][5].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[21][5].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[21][5].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[21][5].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[21][5].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[21][5].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[21][5].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[21][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[21][5].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[21][6].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[21][6].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[21][6].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[21][6].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[21][6].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[21][6].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[21][6].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[21][6].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[21][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[21][6].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[21][7].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[21][7].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[21][7].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[21][7].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[21][7].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[21][7].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[21][7].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[21][7].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[21][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[21][7].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[21][8].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[21][8].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[21][8].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[21][8].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[21][8].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[21][8].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[21][8].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[21][8].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[21][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[21][8].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[21][9].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[21][9].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[21][9].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[21][9].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[21][9].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[21][9].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[21][9].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[21][9].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[21][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[21][9].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[21][10].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[21][10].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[21][10].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[21][10].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[21][10].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[21][10].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[21][10].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[21][10].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[21][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[21][10].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[21][11].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[21][11].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[21][11].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[21][11].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[21][11].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[21][11].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[21][11].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[21][11].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[21][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[21][11].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[21][12].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[21][12].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[21][12].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[21][12].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[21][12].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[21][12].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[21][12].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[21][12].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[21][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[21][12].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[21][13].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[21][13].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[21][13].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[21][13].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[21][13].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[21][13].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[21][13].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[21][13].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[21][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[21][13].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[21][14].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[21][14].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[21][14].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[21][14].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[21][14].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[21][14].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[21][14].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[21][14].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[21][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[21][14].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[21][15].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[21][15].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[21][15].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[21][15].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[21][15].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[21][15].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[21][15].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[21][15].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[21][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[21][15].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[21][16].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[21][16].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[21][16].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[21][16].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[21][16].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[21][16].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[21][16].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[21][16].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[21][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[21][16].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[21][17].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[21][17].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[21][17].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[21][17].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[21][17].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[21][17].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[21][17].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[21][17].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[21][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[21][17].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[21][18].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[21][18].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[21][18].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[21][18].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[21][18].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[21][18].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[21][18].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[21][18].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[21][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[21][18].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[21][19].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[21][19].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[21][19].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[21][19].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[21][19].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[21][19].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[21][19].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[21][19].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[21][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[21][19].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[21][20].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[21][20].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[21][20].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[21][20].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[21][20].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[21][20].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[21][20].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[21][20].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[21][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[21][20].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[21][21].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[21][21].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[21][21].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[21][21].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[21][21].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[21][21].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[21][21].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[21][21].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[21][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[21][21].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[21][22].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[21][22].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[21][22].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[21][22].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[21][22].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[21][22].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[21][22].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[21][22].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[21][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[21][22].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[21][23].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[21][23].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[21][23].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[21][23].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[21][23].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[21][23].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[21][23].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[21][23].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[21][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[21][23].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[21][24].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[21][24].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[21][24].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[21][24].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[21][24].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[21][24].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[21][24].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[21][24].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[21][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[21][24].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[21][25].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[21][25].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[21][25].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[21][25].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[21][25].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[21][25].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[21][25].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[21][25].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[21][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[21][25].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[21][26].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[21][26].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[21][26].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[21][26].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[21][26].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[21][26].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[21][26].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[21][26].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[21][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[21][26].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[21][27].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[21][27].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[21][27].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[21][27].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[21][27].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[21][27].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[21][27].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[21][27].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[21][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[21][27].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[21][28].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[21][28].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[21][28].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[21][28].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[21][28].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[21][28].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[21][28].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[21][28].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[21][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[21][28].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[21][29].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[21][29].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[21][29].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[21][29].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[21][29].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[21][29].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[21][29].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[21][29].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[21][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[21][29].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[21][30].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[21][30].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[21][30].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[21][30].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[21][30].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[21][30].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[21][30].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[21][30].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[21][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[21][30].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[21][31].dma__memc__write_valid      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[21][31].dma__memc__write_address    = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[21][31].dma__memc__write_data       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[21][31].dma__memc__read_valid       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[21][31].dma__memc__read_address     = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[21][31].dma__memc__read_pause       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[21][31].memc__dma__write_ready      = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[21][31].memc__dma__read_data        = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[21][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[21][31].memc__dma__read_ready       = pe_array_inst.pe_inst[21].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 22
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[22][0].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[22][0].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[22][0].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[22][0].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[22][0].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[22][0].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[22][0].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[22][0].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[22][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[22][0].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[22][1].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[22][1].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[22][1].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[22][1].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[22][1].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[22][1].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[22][1].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[22][1].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[22][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[22][1].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[22][2].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[22][2].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[22][2].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[22][2].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[22][2].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[22][2].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[22][2].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[22][2].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[22][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[22][2].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[22][3].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[22][3].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[22][3].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[22][3].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[22][3].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[22][3].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[22][3].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[22][3].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[22][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[22][3].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[22][4].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[22][4].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[22][4].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[22][4].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[22][4].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[22][4].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[22][4].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[22][4].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[22][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[22][4].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[22][5].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[22][5].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[22][5].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[22][5].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[22][5].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[22][5].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[22][5].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[22][5].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[22][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[22][5].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[22][6].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[22][6].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[22][6].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[22][6].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[22][6].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[22][6].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[22][6].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[22][6].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[22][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[22][6].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[22][7].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[22][7].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[22][7].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[22][7].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[22][7].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[22][7].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[22][7].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[22][7].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[22][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[22][7].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[22][8].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[22][8].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[22][8].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[22][8].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[22][8].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[22][8].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[22][8].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[22][8].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[22][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[22][8].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[22][9].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[22][9].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[22][9].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[22][9].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[22][9].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[22][9].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[22][9].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[22][9].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[22][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[22][9].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[22][10].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[22][10].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[22][10].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[22][10].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[22][10].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[22][10].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[22][10].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[22][10].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[22][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[22][10].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[22][11].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[22][11].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[22][11].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[22][11].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[22][11].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[22][11].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[22][11].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[22][11].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[22][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[22][11].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[22][12].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[22][12].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[22][12].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[22][12].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[22][12].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[22][12].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[22][12].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[22][12].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[22][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[22][12].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[22][13].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[22][13].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[22][13].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[22][13].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[22][13].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[22][13].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[22][13].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[22][13].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[22][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[22][13].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[22][14].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[22][14].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[22][14].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[22][14].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[22][14].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[22][14].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[22][14].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[22][14].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[22][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[22][14].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[22][15].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[22][15].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[22][15].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[22][15].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[22][15].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[22][15].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[22][15].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[22][15].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[22][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[22][15].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[22][16].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[22][16].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[22][16].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[22][16].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[22][16].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[22][16].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[22][16].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[22][16].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[22][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[22][16].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[22][17].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[22][17].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[22][17].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[22][17].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[22][17].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[22][17].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[22][17].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[22][17].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[22][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[22][17].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[22][18].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[22][18].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[22][18].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[22][18].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[22][18].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[22][18].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[22][18].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[22][18].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[22][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[22][18].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[22][19].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[22][19].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[22][19].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[22][19].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[22][19].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[22][19].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[22][19].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[22][19].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[22][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[22][19].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[22][20].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[22][20].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[22][20].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[22][20].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[22][20].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[22][20].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[22][20].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[22][20].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[22][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[22][20].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[22][21].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[22][21].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[22][21].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[22][21].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[22][21].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[22][21].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[22][21].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[22][21].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[22][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[22][21].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[22][22].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[22][22].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[22][22].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[22][22].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[22][22].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[22][22].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[22][22].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[22][22].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[22][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[22][22].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[22][23].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[22][23].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[22][23].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[22][23].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[22][23].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[22][23].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[22][23].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[22][23].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[22][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[22][23].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[22][24].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[22][24].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[22][24].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[22][24].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[22][24].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[22][24].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[22][24].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[22][24].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[22][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[22][24].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[22][25].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[22][25].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[22][25].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[22][25].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[22][25].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[22][25].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[22][25].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[22][25].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[22][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[22][25].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[22][26].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[22][26].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[22][26].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[22][26].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[22][26].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[22][26].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[22][26].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[22][26].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[22][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[22][26].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[22][27].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[22][27].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[22][27].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[22][27].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[22][27].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[22][27].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[22][27].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[22][27].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[22][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[22][27].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[22][28].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[22][28].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[22][28].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[22][28].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[22][28].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[22][28].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[22][28].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[22][28].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[22][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[22][28].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[22][29].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[22][29].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[22][29].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[22][29].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[22][29].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[22][29].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[22][29].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[22][29].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[22][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[22][29].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[22][30].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[22][30].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[22][30].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[22][30].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[22][30].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[22][30].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[22][30].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[22][30].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[22][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[22][30].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[22][31].dma__memc__write_valid      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[22][31].dma__memc__write_address    = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[22][31].dma__memc__write_data       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[22][31].dma__memc__read_valid       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[22][31].dma__memc__read_address     = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[22][31].dma__memc__read_pause       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[22][31].memc__dma__write_ready      = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[22][31].memc__dma__read_data        = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[22][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[22][31].memc__dma__read_ready       = pe_array_inst.pe_inst[22].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 23
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[23][0].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[23][0].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[23][0].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[23][0].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[23][0].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[23][0].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[23][0].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[23][0].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[23][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[23][0].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[23][1].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[23][1].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[23][1].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[23][1].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[23][1].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[23][1].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[23][1].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[23][1].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[23][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[23][1].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[23][2].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[23][2].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[23][2].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[23][2].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[23][2].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[23][2].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[23][2].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[23][2].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[23][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[23][2].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[23][3].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[23][3].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[23][3].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[23][3].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[23][3].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[23][3].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[23][3].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[23][3].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[23][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[23][3].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[23][4].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[23][4].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[23][4].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[23][4].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[23][4].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[23][4].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[23][4].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[23][4].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[23][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[23][4].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[23][5].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[23][5].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[23][5].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[23][5].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[23][5].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[23][5].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[23][5].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[23][5].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[23][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[23][5].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[23][6].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[23][6].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[23][6].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[23][6].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[23][6].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[23][6].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[23][6].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[23][6].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[23][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[23][6].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[23][7].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[23][7].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[23][7].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[23][7].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[23][7].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[23][7].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[23][7].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[23][7].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[23][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[23][7].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[23][8].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[23][8].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[23][8].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[23][8].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[23][8].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[23][8].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[23][8].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[23][8].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[23][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[23][8].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[23][9].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[23][9].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[23][9].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[23][9].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[23][9].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[23][9].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[23][9].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[23][9].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[23][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[23][9].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[23][10].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[23][10].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[23][10].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[23][10].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[23][10].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[23][10].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[23][10].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[23][10].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[23][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[23][10].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[23][11].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[23][11].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[23][11].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[23][11].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[23][11].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[23][11].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[23][11].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[23][11].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[23][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[23][11].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[23][12].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[23][12].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[23][12].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[23][12].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[23][12].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[23][12].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[23][12].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[23][12].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[23][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[23][12].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[23][13].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[23][13].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[23][13].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[23][13].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[23][13].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[23][13].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[23][13].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[23][13].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[23][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[23][13].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[23][14].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[23][14].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[23][14].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[23][14].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[23][14].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[23][14].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[23][14].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[23][14].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[23][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[23][14].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[23][15].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[23][15].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[23][15].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[23][15].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[23][15].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[23][15].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[23][15].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[23][15].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[23][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[23][15].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[23][16].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[23][16].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[23][16].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[23][16].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[23][16].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[23][16].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[23][16].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[23][16].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[23][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[23][16].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[23][17].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[23][17].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[23][17].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[23][17].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[23][17].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[23][17].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[23][17].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[23][17].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[23][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[23][17].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[23][18].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[23][18].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[23][18].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[23][18].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[23][18].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[23][18].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[23][18].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[23][18].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[23][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[23][18].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[23][19].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[23][19].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[23][19].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[23][19].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[23][19].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[23][19].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[23][19].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[23][19].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[23][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[23][19].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[23][20].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[23][20].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[23][20].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[23][20].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[23][20].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[23][20].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[23][20].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[23][20].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[23][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[23][20].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[23][21].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[23][21].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[23][21].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[23][21].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[23][21].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[23][21].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[23][21].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[23][21].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[23][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[23][21].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[23][22].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[23][22].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[23][22].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[23][22].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[23][22].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[23][22].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[23][22].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[23][22].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[23][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[23][22].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[23][23].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[23][23].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[23][23].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[23][23].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[23][23].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[23][23].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[23][23].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[23][23].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[23][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[23][23].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[23][24].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[23][24].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[23][24].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[23][24].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[23][24].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[23][24].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[23][24].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[23][24].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[23][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[23][24].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[23][25].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[23][25].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[23][25].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[23][25].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[23][25].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[23][25].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[23][25].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[23][25].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[23][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[23][25].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[23][26].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[23][26].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[23][26].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[23][26].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[23][26].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[23][26].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[23][26].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[23][26].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[23][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[23][26].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[23][27].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[23][27].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[23][27].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[23][27].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[23][27].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[23][27].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[23][27].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[23][27].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[23][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[23][27].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[23][28].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[23][28].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[23][28].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[23][28].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[23][28].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[23][28].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[23][28].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[23][28].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[23][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[23][28].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[23][29].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[23][29].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[23][29].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[23][29].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[23][29].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[23][29].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[23][29].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[23][29].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[23][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[23][29].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[23][30].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[23][30].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[23][30].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[23][30].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[23][30].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[23][30].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[23][30].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[23][30].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[23][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[23][30].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[23][31].dma__memc__write_valid      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[23][31].dma__memc__write_address    = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[23][31].dma__memc__write_data       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[23][31].dma__memc__read_valid       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[23][31].dma__memc__read_address     = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[23][31].dma__memc__read_pause       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[23][31].memc__dma__write_ready      = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[23][31].memc__dma__read_data        = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[23][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[23][31].memc__dma__read_ready       = pe_array_inst.pe_inst[23].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 24
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[24][0].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[24][0].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[24][0].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[24][0].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[24][0].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[24][0].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[24][0].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[24][0].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[24][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[24][0].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[24][1].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[24][1].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[24][1].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[24][1].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[24][1].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[24][1].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[24][1].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[24][1].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[24][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[24][1].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[24][2].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[24][2].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[24][2].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[24][2].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[24][2].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[24][2].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[24][2].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[24][2].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[24][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[24][2].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[24][3].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[24][3].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[24][3].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[24][3].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[24][3].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[24][3].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[24][3].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[24][3].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[24][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[24][3].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[24][4].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[24][4].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[24][4].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[24][4].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[24][4].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[24][4].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[24][4].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[24][4].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[24][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[24][4].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[24][5].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[24][5].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[24][5].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[24][5].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[24][5].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[24][5].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[24][5].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[24][5].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[24][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[24][5].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[24][6].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[24][6].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[24][6].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[24][6].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[24][6].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[24][6].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[24][6].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[24][6].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[24][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[24][6].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[24][7].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[24][7].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[24][7].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[24][7].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[24][7].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[24][7].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[24][7].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[24][7].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[24][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[24][7].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[24][8].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[24][8].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[24][8].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[24][8].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[24][8].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[24][8].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[24][8].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[24][8].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[24][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[24][8].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[24][9].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[24][9].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[24][9].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[24][9].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[24][9].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[24][9].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[24][9].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[24][9].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[24][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[24][9].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[24][10].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[24][10].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[24][10].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[24][10].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[24][10].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[24][10].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[24][10].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[24][10].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[24][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[24][10].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[24][11].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[24][11].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[24][11].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[24][11].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[24][11].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[24][11].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[24][11].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[24][11].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[24][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[24][11].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[24][12].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[24][12].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[24][12].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[24][12].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[24][12].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[24][12].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[24][12].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[24][12].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[24][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[24][12].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[24][13].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[24][13].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[24][13].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[24][13].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[24][13].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[24][13].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[24][13].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[24][13].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[24][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[24][13].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[24][14].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[24][14].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[24][14].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[24][14].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[24][14].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[24][14].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[24][14].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[24][14].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[24][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[24][14].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[24][15].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[24][15].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[24][15].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[24][15].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[24][15].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[24][15].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[24][15].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[24][15].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[24][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[24][15].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[24][16].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[24][16].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[24][16].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[24][16].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[24][16].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[24][16].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[24][16].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[24][16].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[24][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[24][16].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[24][17].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[24][17].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[24][17].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[24][17].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[24][17].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[24][17].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[24][17].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[24][17].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[24][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[24][17].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[24][18].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[24][18].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[24][18].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[24][18].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[24][18].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[24][18].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[24][18].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[24][18].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[24][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[24][18].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[24][19].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[24][19].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[24][19].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[24][19].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[24][19].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[24][19].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[24][19].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[24][19].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[24][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[24][19].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[24][20].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[24][20].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[24][20].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[24][20].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[24][20].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[24][20].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[24][20].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[24][20].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[24][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[24][20].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[24][21].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[24][21].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[24][21].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[24][21].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[24][21].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[24][21].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[24][21].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[24][21].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[24][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[24][21].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[24][22].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[24][22].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[24][22].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[24][22].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[24][22].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[24][22].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[24][22].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[24][22].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[24][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[24][22].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[24][23].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[24][23].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[24][23].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[24][23].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[24][23].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[24][23].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[24][23].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[24][23].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[24][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[24][23].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[24][24].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[24][24].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[24][24].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[24][24].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[24][24].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[24][24].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[24][24].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[24][24].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[24][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[24][24].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[24][25].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[24][25].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[24][25].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[24][25].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[24][25].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[24][25].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[24][25].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[24][25].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[24][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[24][25].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[24][26].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[24][26].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[24][26].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[24][26].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[24][26].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[24][26].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[24][26].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[24][26].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[24][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[24][26].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[24][27].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[24][27].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[24][27].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[24][27].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[24][27].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[24][27].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[24][27].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[24][27].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[24][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[24][27].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[24][28].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[24][28].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[24][28].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[24][28].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[24][28].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[24][28].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[24][28].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[24][28].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[24][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[24][28].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[24][29].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[24][29].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[24][29].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[24][29].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[24][29].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[24][29].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[24][29].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[24][29].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[24][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[24][29].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[24][30].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[24][30].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[24][30].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[24][30].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[24][30].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[24][30].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[24][30].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[24][30].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[24][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[24][30].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[24][31].dma__memc__write_valid      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[24][31].dma__memc__write_address    = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[24][31].dma__memc__write_data       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[24][31].dma__memc__read_valid       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[24][31].dma__memc__read_address     = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[24][31].dma__memc__read_pause       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[24][31].memc__dma__write_ready      = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[24][31].memc__dma__read_data        = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[24][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[24][31].memc__dma__read_ready       = pe_array_inst.pe_inst[24].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 25
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[25][0].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[25][0].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[25][0].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[25][0].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[25][0].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[25][0].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[25][0].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[25][0].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[25][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[25][0].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[25][1].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[25][1].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[25][1].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[25][1].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[25][1].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[25][1].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[25][1].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[25][1].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[25][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[25][1].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[25][2].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[25][2].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[25][2].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[25][2].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[25][2].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[25][2].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[25][2].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[25][2].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[25][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[25][2].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[25][3].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[25][3].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[25][3].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[25][3].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[25][3].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[25][3].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[25][3].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[25][3].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[25][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[25][3].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[25][4].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[25][4].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[25][4].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[25][4].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[25][4].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[25][4].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[25][4].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[25][4].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[25][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[25][4].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[25][5].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[25][5].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[25][5].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[25][5].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[25][5].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[25][5].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[25][5].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[25][5].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[25][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[25][5].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[25][6].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[25][6].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[25][6].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[25][6].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[25][6].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[25][6].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[25][6].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[25][6].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[25][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[25][6].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[25][7].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[25][7].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[25][7].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[25][7].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[25][7].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[25][7].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[25][7].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[25][7].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[25][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[25][7].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[25][8].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[25][8].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[25][8].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[25][8].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[25][8].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[25][8].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[25][8].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[25][8].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[25][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[25][8].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[25][9].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[25][9].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[25][9].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[25][9].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[25][9].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[25][9].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[25][9].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[25][9].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[25][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[25][9].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[25][10].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[25][10].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[25][10].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[25][10].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[25][10].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[25][10].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[25][10].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[25][10].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[25][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[25][10].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[25][11].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[25][11].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[25][11].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[25][11].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[25][11].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[25][11].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[25][11].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[25][11].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[25][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[25][11].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[25][12].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[25][12].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[25][12].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[25][12].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[25][12].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[25][12].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[25][12].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[25][12].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[25][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[25][12].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[25][13].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[25][13].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[25][13].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[25][13].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[25][13].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[25][13].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[25][13].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[25][13].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[25][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[25][13].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[25][14].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[25][14].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[25][14].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[25][14].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[25][14].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[25][14].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[25][14].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[25][14].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[25][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[25][14].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[25][15].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[25][15].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[25][15].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[25][15].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[25][15].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[25][15].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[25][15].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[25][15].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[25][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[25][15].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[25][16].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[25][16].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[25][16].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[25][16].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[25][16].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[25][16].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[25][16].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[25][16].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[25][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[25][16].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[25][17].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[25][17].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[25][17].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[25][17].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[25][17].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[25][17].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[25][17].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[25][17].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[25][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[25][17].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[25][18].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[25][18].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[25][18].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[25][18].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[25][18].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[25][18].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[25][18].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[25][18].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[25][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[25][18].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[25][19].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[25][19].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[25][19].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[25][19].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[25][19].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[25][19].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[25][19].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[25][19].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[25][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[25][19].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[25][20].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[25][20].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[25][20].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[25][20].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[25][20].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[25][20].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[25][20].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[25][20].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[25][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[25][20].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[25][21].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[25][21].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[25][21].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[25][21].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[25][21].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[25][21].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[25][21].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[25][21].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[25][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[25][21].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[25][22].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[25][22].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[25][22].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[25][22].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[25][22].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[25][22].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[25][22].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[25][22].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[25][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[25][22].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[25][23].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[25][23].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[25][23].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[25][23].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[25][23].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[25][23].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[25][23].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[25][23].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[25][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[25][23].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[25][24].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[25][24].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[25][24].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[25][24].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[25][24].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[25][24].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[25][24].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[25][24].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[25][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[25][24].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[25][25].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[25][25].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[25][25].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[25][25].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[25][25].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[25][25].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[25][25].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[25][25].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[25][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[25][25].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[25][26].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[25][26].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[25][26].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[25][26].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[25][26].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[25][26].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[25][26].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[25][26].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[25][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[25][26].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[25][27].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[25][27].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[25][27].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[25][27].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[25][27].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[25][27].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[25][27].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[25][27].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[25][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[25][27].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[25][28].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[25][28].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[25][28].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[25][28].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[25][28].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[25][28].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[25][28].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[25][28].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[25][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[25][28].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[25][29].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[25][29].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[25][29].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[25][29].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[25][29].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[25][29].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[25][29].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[25][29].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[25][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[25][29].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[25][30].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[25][30].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[25][30].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[25][30].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[25][30].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[25][30].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[25][30].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[25][30].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[25][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[25][30].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[25][31].dma__memc__write_valid      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[25][31].dma__memc__write_address    = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[25][31].dma__memc__write_data       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[25][31].dma__memc__read_valid       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[25][31].dma__memc__read_address     = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[25][31].dma__memc__read_pause       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[25][31].memc__dma__write_ready      = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[25][31].memc__dma__read_data        = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[25][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[25][31].memc__dma__read_ready       = pe_array_inst.pe_inst[25].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 26
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[26][0].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[26][0].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[26][0].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[26][0].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[26][0].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[26][0].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[26][0].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[26][0].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[26][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[26][0].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[26][1].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[26][1].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[26][1].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[26][1].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[26][1].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[26][1].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[26][1].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[26][1].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[26][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[26][1].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[26][2].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[26][2].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[26][2].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[26][2].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[26][2].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[26][2].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[26][2].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[26][2].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[26][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[26][2].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[26][3].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[26][3].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[26][3].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[26][3].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[26][3].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[26][3].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[26][3].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[26][3].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[26][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[26][3].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[26][4].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[26][4].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[26][4].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[26][4].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[26][4].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[26][4].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[26][4].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[26][4].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[26][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[26][4].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[26][5].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[26][5].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[26][5].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[26][5].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[26][5].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[26][5].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[26][5].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[26][5].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[26][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[26][5].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[26][6].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[26][6].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[26][6].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[26][6].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[26][6].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[26][6].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[26][6].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[26][6].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[26][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[26][6].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[26][7].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[26][7].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[26][7].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[26][7].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[26][7].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[26][7].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[26][7].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[26][7].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[26][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[26][7].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[26][8].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[26][8].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[26][8].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[26][8].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[26][8].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[26][8].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[26][8].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[26][8].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[26][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[26][8].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[26][9].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[26][9].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[26][9].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[26][9].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[26][9].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[26][9].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[26][9].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[26][9].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[26][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[26][9].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[26][10].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[26][10].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[26][10].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[26][10].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[26][10].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[26][10].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[26][10].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[26][10].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[26][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[26][10].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[26][11].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[26][11].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[26][11].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[26][11].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[26][11].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[26][11].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[26][11].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[26][11].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[26][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[26][11].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[26][12].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[26][12].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[26][12].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[26][12].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[26][12].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[26][12].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[26][12].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[26][12].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[26][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[26][12].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[26][13].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[26][13].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[26][13].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[26][13].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[26][13].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[26][13].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[26][13].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[26][13].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[26][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[26][13].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[26][14].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[26][14].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[26][14].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[26][14].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[26][14].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[26][14].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[26][14].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[26][14].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[26][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[26][14].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[26][15].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[26][15].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[26][15].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[26][15].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[26][15].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[26][15].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[26][15].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[26][15].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[26][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[26][15].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[26][16].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[26][16].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[26][16].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[26][16].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[26][16].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[26][16].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[26][16].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[26][16].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[26][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[26][16].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[26][17].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[26][17].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[26][17].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[26][17].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[26][17].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[26][17].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[26][17].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[26][17].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[26][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[26][17].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[26][18].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[26][18].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[26][18].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[26][18].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[26][18].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[26][18].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[26][18].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[26][18].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[26][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[26][18].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[26][19].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[26][19].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[26][19].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[26][19].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[26][19].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[26][19].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[26][19].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[26][19].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[26][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[26][19].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[26][20].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[26][20].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[26][20].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[26][20].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[26][20].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[26][20].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[26][20].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[26][20].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[26][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[26][20].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[26][21].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[26][21].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[26][21].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[26][21].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[26][21].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[26][21].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[26][21].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[26][21].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[26][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[26][21].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[26][22].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[26][22].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[26][22].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[26][22].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[26][22].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[26][22].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[26][22].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[26][22].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[26][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[26][22].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[26][23].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[26][23].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[26][23].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[26][23].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[26][23].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[26][23].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[26][23].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[26][23].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[26][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[26][23].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[26][24].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[26][24].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[26][24].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[26][24].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[26][24].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[26][24].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[26][24].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[26][24].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[26][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[26][24].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[26][25].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[26][25].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[26][25].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[26][25].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[26][25].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[26][25].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[26][25].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[26][25].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[26][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[26][25].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[26][26].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[26][26].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[26][26].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[26][26].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[26][26].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[26][26].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[26][26].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[26][26].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[26][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[26][26].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[26][27].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[26][27].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[26][27].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[26][27].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[26][27].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[26][27].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[26][27].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[26][27].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[26][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[26][27].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[26][28].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[26][28].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[26][28].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[26][28].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[26][28].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[26][28].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[26][28].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[26][28].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[26][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[26][28].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[26][29].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[26][29].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[26][29].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[26][29].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[26][29].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[26][29].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[26][29].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[26][29].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[26][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[26][29].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[26][30].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[26][30].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[26][30].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[26][30].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[26][30].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[26][30].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[26][30].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[26][30].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[26][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[26][30].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[26][31].dma__memc__write_valid      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[26][31].dma__memc__write_address    = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[26][31].dma__memc__write_data       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[26][31].dma__memc__read_valid       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[26][31].dma__memc__read_address     = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[26][31].dma__memc__read_pause       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[26][31].memc__dma__write_ready      = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[26][31].memc__dma__read_data        = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[26][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[26][31].memc__dma__read_ready       = pe_array_inst.pe_inst[26].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 27
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[27][0].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[27][0].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[27][0].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[27][0].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[27][0].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[27][0].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[27][0].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[27][0].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[27][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[27][0].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[27][1].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[27][1].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[27][1].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[27][1].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[27][1].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[27][1].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[27][1].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[27][1].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[27][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[27][1].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[27][2].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[27][2].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[27][2].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[27][2].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[27][2].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[27][2].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[27][2].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[27][2].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[27][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[27][2].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[27][3].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[27][3].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[27][3].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[27][3].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[27][3].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[27][3].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[27][3].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[27][3].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[27][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[27][3].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[27][4].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[27][4].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[27][4].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[27][4].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[27][4].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[27][4].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[27][4].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[27][4].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[27][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[27][4].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[27][5].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[27][5].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[27][5].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[27][5].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[27][5].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[27][5].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[27][5].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[27][5].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[27][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[27][5].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[27][6].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[27][6].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[27][6].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[27][6].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[27][6].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[27][6].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[27][6].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[27][6].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[27][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[27][6].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[27][7].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[27][7].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[27][7].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[27][7].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[27][7].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[27][7].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[27][7].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[27][7].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[27][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[27][7].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[27][8].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[27][8].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[27][8].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[27][8].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[27][8].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[27][8].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[27][8].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[27][8].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[27][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[27][8].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[27][9].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[27][9].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[27][9].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[27][9].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[27][9].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[27][9].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[27][9].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[27][9].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[27][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[27][9].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[27][10].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[27][10].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[27][10].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[27][10].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[27][10].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[27][10].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[27][10].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[27][10].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[27][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[27][10].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[27][11].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[27][11].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[27][11].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[27][11].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[27][11].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[27][11].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[27][11].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[27][11].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[27][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[27][11].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[27][12].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[27][12].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[27][12].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[27][12].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[27][12].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[27][12].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[27][12].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[27][12].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[27][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[27][12].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[27][13].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[27][13].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[27][13].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[27][13].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[27][13].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[27][13].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[27][13].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[27][13].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[27][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[27][13].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[27][14].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[27][14].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[27][14].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[27][14].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[27][14].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[27][14].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[27][14].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[27][14].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[27][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[27][14].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[27][15].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[27][15].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[27][15].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[27][15].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[27][15].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[27][15].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[27][15].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[27][15].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[27][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[27][15].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[27][16].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[27][16].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[27][16].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[27][16].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[27][16].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[27][16].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[27][16].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[27][16].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[27][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[27][16].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[27][17].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[27][17].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[27][17].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[27][17].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[27][17].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[27][17].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[27][17].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[27][17].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[27][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[27][17].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[27][18].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[27][18].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[27][18].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[27][18].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[27][18].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[27][18].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[27][18].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[27][18].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[27][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[27][18].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[27][19].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[27][19].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[27][19].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[27][19].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[27][19].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[27][19].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[27][19].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[27][19].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[27][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[27][19].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[27][20].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[27][20].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[27][20].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[27][20].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[27][20].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[27][20].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[27][20].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[27][20].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[27][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[27][20].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[27][21].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[27][21].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[27][21].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[27][21].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[27][21].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[27][21].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[27][21].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[27][21].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[27][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[27][21].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[27][22].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[27][22].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[27][22].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[27][22].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[27][22].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[27][22].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[27][22].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[27][22].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[27][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[27][22].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[27][23].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[27][23].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[27][23].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[27][23].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[27][23].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[27][23].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[27][23].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[27][23].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[27][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[27][23].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[27][24].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[27][24].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[27][24].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[27][24].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[27][24].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[27][24].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[27][24].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[27][24].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[27][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[27][24].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[27][25].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[27][25].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[27][25].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[27][25].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[27][25].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[27][25].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[27][25].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[27][25].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[27][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[27][25].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[27][26].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[27][26].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[27][26].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[27][26].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[27][26].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[27][26].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[27][26].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[27][26].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[27][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[27][26].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[27][27].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[27][27].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[27][27].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[27][27].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[27][27].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[27][27].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[27][27].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[27][27].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[27][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[27][27].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[27][28].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[27][28].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[27][28].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[27][28].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[27][28].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[27][28].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[27][28].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[27][28].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[27][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[27][28].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[27][29].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[27][29].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[27][29].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[27][29].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[27][29].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[27][29].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[27][29].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[27][29].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[27][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[27][29].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[27][30].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[27][30].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[27][30].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[27][30].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[27][30].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[27][30].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[27][30].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[27][30].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[27][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[27][30].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[27][31].dma__memc__write_valid      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[27][31].dma__memc__write_address    = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[27][31].dma__memc__write_data       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[27][31].dma__memc__read_valid       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[27][31].dma__memc__read_address     = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[27][31].dma__memc__read_pause       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[27][31].memc__dma__write_ready      = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[27][31].memc__dma__read_data        = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[27][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[27][31].memc__dma__read_ready       = pe_array_inst.pe_inst[27].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 28
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[28][0].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[28][0].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[28][0].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[28][0].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[28][0].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[28][0].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[28][0].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[28][0].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[28][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[28][0].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[28][1].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[28][1].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[28][1].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[28][1].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[28][1].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[28][1].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[28][1].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[28][1].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[28][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[28][1].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[28][2].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[28][2].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[28][2].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[28][2].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[28][2].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[28][2].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[28][2].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[28][2].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[28][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[28][2].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[28][3].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[28][3].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[28][3].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[28][3].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[28][3].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[28][3].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[28][3].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[28][3].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[28][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[28][3].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[28][4].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[28][4].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[28][4].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[28][4].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[28][4].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[28][4].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[28][4].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[28][4].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[28][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[28][4].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[28][5].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[28][5].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[28][5].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[28][5].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[28][5].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[28][5].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[28][5].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[28][5].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[28][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[28][5].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[28][6].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[28][6].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[28][6].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[28][6].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[28][6].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[28][6].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[28][6].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[28][6].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[28][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[28][6].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[28][7].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[28][7].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[28][7].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[28][7].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[28][7].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[28][7].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[28][7].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[28][7].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[28][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[28][7].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[28][8].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[28][8].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[28][8].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[28][8].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[28][8].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[28][8].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[28][8].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[28][8].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[28][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[28][8].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[28][9].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[28][9].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[28][9].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[28][9].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[28][9].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[28][9].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[28][9].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[28][9].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[28][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[28][9].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[28][10].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[28][10].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[28][10].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[28][10].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[28][10].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[28][10].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[28][10].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[28][10].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[28][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[28][10].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[28][11].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[28][11].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[28][11].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[28][11].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[28][11].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[28][11].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[28][11].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[28][11].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[28][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[28][11].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[28][12].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[28][12].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[28][12].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[28][12].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[28][12].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[28][12].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[28][12].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[28][12].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[28][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[28][12].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[28][13].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[28][13].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[28][13].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[28][13].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[28][13].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[28][13].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[28][13].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[28][13].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[28][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[28][13].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[28][14].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[28][14].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[28][14].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[28][14].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[28][14].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[28][14].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[28][14].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[28][14].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[28][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[28][14].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[28][15].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[28][15].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[28][15].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[28][15].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[28][15].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[28][15].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[28][15].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[28][15].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[28][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[28][15].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[28][16].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[28][16].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[28][16].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[28][16].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[28][16].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[28][16].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[28][16].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[28][16].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[28][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[28][16].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[28][17].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[28][17].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[28][17].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[28][17].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[28][17].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[28][17].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[28][17].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[28][17].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[28][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[28][17].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[28][18].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[28][18].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[28][18].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[28][18].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[28][18].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[28][18].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[28][18].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[28][18].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[28][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[28][18].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[28][19].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[28][19].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[28][19].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[28][19].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[28][19].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[28][19].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[28][19].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[28][19].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[28][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[28][19].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[28][20].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[28][20].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[28][20].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[28][20].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[28][20].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[28][20].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[28][20].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[28][20].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[28][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[28][20].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[28][21].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[28][21].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[28][21].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[28][21].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[28][21].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[28][21].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[28][21].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[28][21].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[28][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[28][21].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[28][22].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[28][22].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[28][22].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[28][22].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[28][22].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[28][22].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[28][22].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[28][22].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[28][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[28][22].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[28][23].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[28][23].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[28][23].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[28][23].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[28][23].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[28][23].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[28][23].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[28][23].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[28][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[28][23].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[28][24].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[28][24].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[28][24].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[28][24].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[28][24].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[28][24].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[28][24].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[28][24].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[28][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[28][24].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[28][25].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[28][25].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[28][25].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[28][25].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[28][25].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[28][25].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[28][25].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[28][25].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[28][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[28][25].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[28][26].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[28][26].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[28][26].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[28][26].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[28][26].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[28][26].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[28][26].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[28][26].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[28][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[28][26].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[28][27].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[28][27].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[28][27].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[28][27].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[28][27].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[28][27].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[28][27].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[28][27].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[28][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[28][27].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[28][28].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[28][28].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[28][28].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[28][28].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[28][28].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[28][28].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[28][28].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[28][28].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[28][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[28][28].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[28][29].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[28][29].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[28][29].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[28][29].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[28][29].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[28][29].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[28][29].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[28][29].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[28][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[28][29].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[28][30].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[28][30].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[28][30].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[28][30].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[28][30].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[28][30].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[28][30].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[28][30].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[28][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[28][30].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[28][31].dma__memc__write_valid      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[28][31].dma__memc__write_address    = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[28][31].dma__memc__write_data       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[28][31].dma__memc__read_valid       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[28][31].dma__memc__read_address     = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[28][31].dma__memc__read_pause       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[28][31].memc__dma__write_ready      = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[28][31].memc__dma__read_data        = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[28][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[28][31].memc__dma__read_ready       = pe_array_inst.pe_inst[28].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 29
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[29][0].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[29][0].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[29][0].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[29][0].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[29][0].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[29][0].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[29][0].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[29][0].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[29][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[29][0].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[29][1].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[29][1].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[29][1].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[29][1].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[29][1].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[29][1].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[29][1].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[29][1].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[29][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[29][1].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[29][2].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[29][2].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[29][2].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[29][2].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[29][2].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[29][2].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[29][2].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[29][2].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[29][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[29][2].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[29][3].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[29][3].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[29][3].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[29][3].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[29][3].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[29][3].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[29][3].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[29][3].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[29][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[29][3].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[29][4].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[29][4].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[29][4].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[29][4].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[29][4].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[29][4].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[29][4].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[29][4].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[29][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[29][4].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[29][5].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[29][5].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[29][5].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[29][5].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[29][5].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[29][5].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[29][5].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[29][5].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[29][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[29][5].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[29][6].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[29][6].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[29][6].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[29][6].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[29][6].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[29][6].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[29][6].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[29][6].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[29][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[29][6].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[29][7].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[29][7].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[29][7].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[29][7].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[29][7].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[29][7].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[29][7].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[29][7].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[29][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[29][7].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[29][8].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[29][8].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[29][8].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[29][8].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[29][8].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[29][8].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[29][8].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[29][8].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[29][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[29][8].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[29][9].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[29][9].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[29][9].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[29][9].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[29][9].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[29][9].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[29][9].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[29][9].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[29][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[29][9].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[29][10].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[29][10].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[29][10].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[29][10].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[29][10].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[29][10].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[29][10].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[29][10].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[29][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[29][10].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[29][11].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[29][11].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[29][11].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[29][11].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[29][11].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[29][11].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[29][11].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[29][11].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[29][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[29][11].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[29][12].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[29][12].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[29][12].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[29][12].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[29][12].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[29][12].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[29][12].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[29][12].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[29][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[29][12].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[29][13].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[29][13].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[29][13].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[29][13].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[29][13].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[29][13].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[29][13].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[29][13].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[29][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[29][13].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[29][14].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[29][14].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[29][14].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[29][14].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[29][14].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[29][14].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[29][14].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[29][14].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[29][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[29][14].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[29][15].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[29][15].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[29][15].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[29][15].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[29][15].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[29][15].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[29][15].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[29][15].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[29][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[29][15].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[29][16].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[29][16].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[29][16].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[29][16].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[29][16].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[29][16].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[29][16].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[29][16].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[29][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[29][16].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[29][17].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[29][17].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[29][17].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[29][17].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[29][17].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[29][17].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[29][17].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[29][17].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[29][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[29][17].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[29][18].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[29][18].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[29][18].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[29][18].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[29][18].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[29][18].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[29][18].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[29][18].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[29][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[29][18].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[29][19].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[29][19].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[29][19].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[29][19].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[29][19].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[29][19].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[29][19].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[29][19].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[29][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[29][19].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[29][20].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[29][20].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[29][20].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[29][20].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[29][20].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[29][20].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[29][20].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[29][20].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[29][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[29][20].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[29][21].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[29][21].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[29][21].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[29][21].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[29][21].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[29][21].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[29][21].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[29][21].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[29][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[29][21].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[29][22].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[29][22].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[29][22].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[29][22].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[29][22].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[29][22].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[29][22].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[29][22].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[29][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[29][22].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[29][23].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[29][23].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[29][23].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[29][23].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[29][23].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[29][23].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[29][23].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[29][23].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[29][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[29][23].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[29][24].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[29][24].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[29][24].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[29][24].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[29][24].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[29][24].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[29][24].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[29][24].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[29][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[29][24].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[29][25].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[29][25].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[29][25].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[29][25].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[29][25].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[29][25].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[29][25].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[29][25].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[29][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[29][25].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[29][26].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[29][26].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[29][26].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[29][26].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[29][26].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[29][26].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[29][26].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[29][26].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[29][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[29][26].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[29][27].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[29][27].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[29][27].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[29][27].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[29][27].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[29][27].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[29][27].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[29][27].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[29][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[29][27].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[29][28].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[29][28].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[29][28].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[29][28].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[29][28].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[29][28].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[29][28].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[29][28].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[29][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[29][28].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[29][29].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[29][29].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[29][29].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[29][29].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[29][29].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[29][29].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[29][29].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[29][29].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[29][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[29][29].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[29][30].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[29][30].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[29][30].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[29][30].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[29][30].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[29][30].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[29][30].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[29][30].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[29][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[29][30].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[29][31].dma__memc__write_valid      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[29][31].dma__memc__write_address    = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[29][31].dma__memc__write_data       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[29][31].dma__memc__read_valid       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[29][31].dma__memc__read_address     = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[29][31].dma__memc__read_pause       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[29][31].memc__dma__write_ready      = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[29][31].memc__dma__read_data        = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[29][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[29][31].memc__dma__read_ready       = pe_array_inst.pe_inst[29].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 30
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[30][0].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[30][0].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[30][0].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[30][0].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[30][0].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[30][0].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[30][0].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[30][0].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[30][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[30][0].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[30][1].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[30][1].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[30][1].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[30][1].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[30][1].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[30][1].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[30][1].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[30][1].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[30][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[30][1].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[30][2].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[30][2].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[30][2].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[30][2].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[30][2].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[30][2].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[30][2].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[30][2].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[30][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[30][2].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[30][3].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[30][3].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[30][3].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[30][3].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[30][3].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[30][3].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[30][3].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[30][3].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[30][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[30][3].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[30][4].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[30][4].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[30][4].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[30][4].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[30][4].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[30][4].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[30][4].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[30][4].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[30][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[30][4].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[30][5].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[30][5].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[30][5].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[30][5].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[30][5].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[30][5].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[30][5].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[30][5].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[30][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[30][5].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[30][6].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[30][6].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[30][6].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[30][6].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[30][6].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[30][6].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[30][6].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[30][6].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[30][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[30][6].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[30][7].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[30][7].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[30][7].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[30][7].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[30][7].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[30][7].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[30][7].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[30][7].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[30][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[30][7].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[30][8].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[30][8].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[30][8].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[30][8].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[30][8].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[30][8].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[30][8].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[30][8].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[30][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[30][8].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[30][9].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[30][9].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[30][9].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[30][9].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[30][9].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[30][9].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[30][9].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[30][9].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[30][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[30][9].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[30][10].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[30][10].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[30][10].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[30][10].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[30][10].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[30][10].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[30][10].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[30][10].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[30][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[30][10].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[30][11].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[30][11].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[30][11].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[30][11].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[30][11].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[30][11].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[30][11].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[30][11].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[30][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[30][11].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[30][12].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[30][12].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[30][12].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[30][12].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[30][12].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[30][12].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[30][12].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[30][12].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[30][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[30][12].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[30][13].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[30][13].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[30][13].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[30][13].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[30][13].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[30][13].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[30][13].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[30][13].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[30][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[30][13].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[30][14].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[30][14].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[30][14].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[30][14].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[30][14].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[30][14].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[30][14].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[30][14].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[30][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[30][14].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[30][15].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[30][15].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[30][15].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[30][15].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[30][15].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[30][15].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[30][15].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[30][15].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[30][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[30][15].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[30][16].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[30][16].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[30][16].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[30][16].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[30][16].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[30][16].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[30][16].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[30][16].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[30][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[30][16].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[30][17].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[30][17].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[30][17].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[30][17].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[30][17].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[30][17].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[30][17].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[30][17].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[30][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[30][17].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[30][18].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[30][18].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[30][18].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[30][18].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[30][18].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[30][18].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[30][18].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[30][18].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[30][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[30][18].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[30][19].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[30][19].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[30][19].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[30][19].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[30][19].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[30][19].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[30][19].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[30][19].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[30][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[30][19].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[30][20].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[30][20].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[30][20].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[30][20].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[30][20].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[30][20].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[30][20].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[30][20].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[30][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[30][20].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[30][21].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[30][21].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[30][21].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[30][21].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[30][21].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[30][21].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[30][21].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[30][21].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[30][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[30][21].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[30][22].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[30][22].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[30][22].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[30][22].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[30][22].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[30][22].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[30][22].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[30][22].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[30][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[30][22].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[30][23].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[30][23].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[30][23].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[30][23].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[30][23].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[30][23].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[30][23].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[30][23].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[30][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[30][23].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[30][24].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[30][24].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[30][24].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[30][24].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[30][24].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[30][24].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[30][24].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[30][24].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[30][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[30][24].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[30][25].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[30][25].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[30][25].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[30][25].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[30][25].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[30][25].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[30][25].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[30][25].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[30][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[30][25].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[30][26].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[30][26].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[30][26].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[30][26].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[30][26].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[30][26].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[30][26].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[30][26].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[30][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[30][26].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[30][27].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[30][27].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[30][27].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[30][27].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[30][27].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[30][27].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[30][27].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[30][27].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[30][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[30][27].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[30][28].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[30][28].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[30][28].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[30][28].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[30][28].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[30][28].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[30][28].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[30][28].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[30][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[30][28].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[30][29].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[30][29].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[30][29].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[30][29].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[30][29].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[30][29].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[30][29].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[30][29].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[30][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[30][29].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[30][30].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[30][30].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[30][30].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[30][30].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[30][30].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[30][30].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[30][30].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[30][30].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[30][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[30][30].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[30][31].dma__memc__write_valid      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[30][31].dma__memc__write_address    = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[30][31].dma__memc__write_data       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[30][31].dma__memc__read_valid       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[30][31].dma__memc__read_address     = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[30][31].dma__memc__read_pause       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[30][31].memc__dma__write_ready      = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[30][31].memc__dma__read_data        = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[30][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[30][31].memc__dma__read_ready       = pe_array_inst.pe_inst[30].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 31
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[31][0].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[31][0].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[31][0].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[31][0].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[31][0].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[31][0].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[31][0].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[31][0].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[31][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[31][0].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[31][1].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[31][1].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[31][1].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[31][1].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[31][1].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[31][1].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[31][1].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[31][1].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[31][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[31][1].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[31][2].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[31][2].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[31][2].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[31][2].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[31][2].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[31][2].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[31][2].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[31][2].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[31][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[31][2].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[31][3].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[31][3].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[31][3].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[31][3].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[31][3].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[31][3].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[31][3].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[31][3].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[31][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[31][3].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[31][4].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[31][4].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[31][4].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[31][4].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[31][4].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[31][4].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[31][4].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[31][4].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[31][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[31][4].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[31][5].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[31][5].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[31][5].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[31][5].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[31][5].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[31][5].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[31][5].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[31][5].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[31][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[31][5].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[31][6].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[31][6].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[31][6].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[31][6].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[31][6].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[31][6].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[31][6].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[31][6].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[31][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[31][6].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[31][7].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[31][7].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[31][7].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[31][7].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[31][7].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[31][7].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[31][7].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[31][7].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[31][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[31][7].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[31][8].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[31][8].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[31][8].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[31][8].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[31][8].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[31][8].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[31][8].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[31][8].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[31][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[31][8].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[31][9].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[31][9].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[31][9].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[31][9].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[31][9].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[31][9].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[31][9].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[31][9].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[31][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[31][9].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[31][10].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[31][10].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[31][10].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[31][10].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[31][10].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[31][10].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[31][10].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[31][10].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[31][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[31][10].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[31][11].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[31][11].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[31][11].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[31][11].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[31][11].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[31][11].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[31][11].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[31][11].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[31][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[31][11].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[31][12].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[31][12].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[31][12].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[31][12].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[31][12].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[31][12].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[31][12].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[31][12].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[31][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[31][12].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[31][13].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[31][13].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[31][13].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[31][13].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[31][13].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[31][13].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[31][13].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[31][13].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[31][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[31][13].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[31][14].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[31][14].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[31][14].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[31][14].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[31][14].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[31][14].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[31][14].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[31][14].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[31][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[31][14].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[31][15].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[31][15].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[31][15].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[31][15].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[31][15].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[31][15].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[31][15].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[31][15].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[31][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[31][15].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[31][16].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[31][16].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[31][16].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[31][16].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[31][16].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[31][16].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[31][16].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[31][16].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[31][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[31][16].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[31][17].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[31][17].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[31][17].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[31][17].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[31][17].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[31][17].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[31][17].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[31][17].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[31][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[31][17].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[31][18].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[31][18].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[31][18].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[31][18].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[31][18].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[31][18].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[31][18].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[31][18].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[31][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[31][18].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[31][19].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[31][19].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[31][19].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[31][19].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[31][19].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[31][19].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[31][19].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[31][19].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[31][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[31][19].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[31][20].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[31][20].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[31][20].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[31][20].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[31][20].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[31][20].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[31][20].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[31][20].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[31][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[31][20].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[31][21].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[31][21].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[31][21].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[31][21].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[31][21].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[31][21].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[31][21].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[31][21].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[31][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[31][21].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[31][22].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[31][22].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[31][22].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[31][22].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[31][22].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[31][22].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[31][22].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[31][22].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[31][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[31][22].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[31][23].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[31][23].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[31][23].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[31][23].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[31][23].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[31][23].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[31][23].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[31][23].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[31][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[31][23].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[31][24].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[31][24].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[31][24].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[31][24].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[31][24].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[31][24].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[31][24].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[31][24].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[31][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[31][24].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[31][25].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[31][25].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[31][25].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[31][25].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[31][25].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[31][25].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[31][25].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[31][25].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[31][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[31][25].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[31][26].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[31][26].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[31][26].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[31][26].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[31][26].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[31][26].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[31][26].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[31][26].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[31][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[31][26].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[31][27].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[31][27].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[31][27].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[31][27].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[31][27].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[31][27].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[31][27].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[31][27].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[31][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[31][27].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[31][28].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[31][28].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[31][28].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[31][28].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[31][28].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[31][28].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[31][28].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[31][28].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[31][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[31][28].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[31][29].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[31][29].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[31][29].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[31][29].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[31][29].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[31][29].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[31][29].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[31][29].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[31][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[31][29].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[31][30].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[31][30].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[31][30].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[31][30].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[31][30].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[31][30].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[31][30].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[31][30].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[31][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[31][30].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[31][31].dma__memc__write_valid      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[31][31].dma__memc__write_address    = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[31][31].dma__memc__write_data       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[31][31].dma__memc__read_valid       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[31][31].dma__memc__read_address     = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[31][31].dma__memc__read_pause       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[31][31].memc__dma__write_ready      = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[31][31].memc__dma__read_data        = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[31][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[31][31].memc__dma__read_ready       = pe_array_inst.pe_inst[31].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 32
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[32][0].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[32][0].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[32][0].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[32][0].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[32][0].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[32][0].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[32][0].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[32][0].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[32][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[32][0].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[32][1].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[32][1].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[32][1].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[32][1].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[32][1].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[32][1].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[32][1].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[32][1].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[32][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[32][1].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[32][2].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[32][2].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[32][2].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[32][2].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[32][2].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[32][2].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[32][2].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[32][2].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[32][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[32][2].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[32][3].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[32][3].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[32][3].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[32][3].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[32][3].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[32][3].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[32][3].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[32][3].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[32][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[32][3].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[32][4].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[32][4].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[32][4].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[32][4].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[32][4].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[32][4].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[32][4].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[32][4].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[32][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[32][4].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[32][5].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[32][5].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[32][5].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[32][5].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[32][5].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[32][5].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[32][5].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[32][5].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[32][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[32][5].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[32][6].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[32][6].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[32][6].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[32][6].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[32][6].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[32][6].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[32][6].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[32][6].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[32][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[32][6].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[32][7].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[32][7].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[32][7].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[32][7].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[32][7].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[32][7].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[32][7].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[32][7].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[32][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[32][7].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[32][8].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[32][8].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[32][8].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[32][8].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[32][8].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[32][8].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[32][8].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[32][8].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[32][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[32][8].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[32][9].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[32][9].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[32][9].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[32][9].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[32][9].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[32][9].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[32][9].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[32][9].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[32][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[32][9].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[32][10].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[32][10].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[32][10].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[32][10].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[32][10].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[32][10].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[32][10].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[32][10].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[32][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[32][10].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[32][11].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[32][11].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[32][11].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[32][11].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[32][11].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[32][11].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[32][11].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[32][11].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[32][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[32][11].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[32][12].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[32][12].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[32][12].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[32][12].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[32][12].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[32][12].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[32][12].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[32][12].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[32][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[32][12].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[32][13].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[32][13].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[32][13].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[32][13].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[32][13].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[32][13].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[32][13].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[32][13].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[32][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[32][13].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[32][14].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[32][14].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[32][14].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[32][14].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[32][14].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[32][14].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[32][14].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[32][14].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[32][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[32][14].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[32][15].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[32][15].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[32][15].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[32][15].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[32][15].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[32][15].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[32][15].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[32][15].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[32][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[32][15].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[32][16].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[32][16].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[32][16].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[32][16].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[32][16].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[32][16].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[32][16].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[32][16].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[32][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[32][16].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[32][17].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[32][17].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[32][17].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[32][17].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[32][17].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[32][17].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[32][17].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[32][17].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[32][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[32][17].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[32][18].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[32][18].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[32][18].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[32][18].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[32][18].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[32][18].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[32][18].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[32][18].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[32][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[32][18].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[32][19].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[32][19].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[32][19].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[32][19].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[32][19].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[32][19].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[32][19].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[32][19].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[32][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[32][19].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[32][20].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[32][20].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[32][20].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[32][20].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[32][20].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[32][20].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[32][20].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[32][20].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[32][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[32][20].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[32][21].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[32][21].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[32][21].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[32][21].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[32][21].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[32][21].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[32][21].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[32][21].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[32][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[32][21].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[32][22].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[32][22].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[32][22].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[32][22].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[32][22].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[32][22].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[32][22].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[32][22].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[32][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[32][22].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[32][23].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[32][23].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[32][23].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[32][23].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[32][23].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[32][23].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[32][23].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[32][23].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[32][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[32][23].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[32][24].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[32][24].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[32][24].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[32][24].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[32][24].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[32][24].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[32][24].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[32][24].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[32][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[32][24].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[32][25].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[32][25].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[32][25].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[32][25].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[32][25].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[32][25].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[32][25].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[32][25].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[32][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[32][25].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[32][26].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[32][26].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[32][26].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[32][26].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[32][26].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[32][26].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[32][26].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[32][26].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[32][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[32][26].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[32][27].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[32][27].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[32][27].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[32][27].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[32][27].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[32][27].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[32][27].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[32][27].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[32][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[32][27].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[32][28].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[32][28].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[32][28].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[32][28].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[32][28].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[32][28].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[32][28].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[32][28].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[32][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[32][28].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[32][29].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[32][29].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[32][29].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[32][29].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[32][29].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[32][29].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[32][29].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[32][29].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[32][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[32][29].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[32][30].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[32][30].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[32][30].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[32][30].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[32][30].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[32][30].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[32][30].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[32][30].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[32][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[32][30].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[32][31].dma__memc__write_valid      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[32][31].dma__memc__write_address    = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[32][31].dma__memc__write_data       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[32][31].dma__memc__read_valid       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[32][31].dma__memc__read_address     = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[32][31].dma__memc__read_pause       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[32][31].memc__dma__write_ready      = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[32][31].memc__dma__read_data        = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[32][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[32][31].memc__dma__read_ready       = pe_array_inst.pe_inst[32].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 33
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[33][0].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[33][0].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[33][0].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[33][0].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[33][0].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[33][0].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[33][0].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[33][0].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[33][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[33][0].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[33][1].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[33][1].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[33][1].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[33][1].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[33][1].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[33][1].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[33][1].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[33][1].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[33][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[33][1].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[33][2].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[33][2].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[33][2].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[33][2].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[33][2].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[33][2].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[33][2].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[33][2].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[33][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[33][2].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[33][3].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[33][3].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[33][3].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[33][3].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[33][3].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[33][3].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[33][3].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[33][3].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[33][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[33][3].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[33][4].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[33][4].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[33][4].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[33][4].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[33][4].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[33][4].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[33][4].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[33][4].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[33][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[33][4].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[33][5].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[33][5].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[33][5].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[33][5].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[33][5].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[33][5].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[33][5].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[33][5].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[33][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[33][5].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[33][6].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[33][6].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[33][6].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[33][6].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[33][6].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[33][6].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[33][6].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[33][6].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[33][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[33][6].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[33][7].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[33][7].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[33][7].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[33][7].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[33][7].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[33][7].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[33][7].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[33][7].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[33][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[33][7].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[33][8].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[33][8].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[33][8].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[33][8].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[33][8].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[33][8].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[33][8].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[33][8].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[33][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[33][8].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[33][9].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[33][9].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[33][9].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[33][9].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[33][9].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[33][9].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[33][9].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[33][9].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[33][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[33][9].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[33][10].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[33][10].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[33][10].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[33][10].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[33][10].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[33][10].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[33][10].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[33][10].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[33][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[33][10].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[33][11].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[33][11].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[33][11].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[33][11].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[33][11].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[33][11].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[33][11].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[33][11].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[33][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[33][11].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[33][12].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[33][12].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[33][12].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[33][12].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[33][12].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[33][12].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[33][12].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[33][12].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[33][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[33][12].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[33][13].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[33][13].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[33][13].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[33][13].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[33][13].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[33][13].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[33][13].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[33][13].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[33][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[33][13].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[33][14].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[33][14].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[33][14].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[33][14].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[33][14].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[33][14].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[33][14].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[33][14].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[33][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[33][14].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[33][15].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[33][15].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[33][15].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[33][15].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[33][15].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[33][15].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[33][15].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[33][15].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[33][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[33][15].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[33][16].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[33][16].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[33][16].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[33][16].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[33][16].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[33][16].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[33][16].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[33][16].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[33][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[33][16].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[33][17].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[33][17].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[33][17].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[33][17].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[33][17].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[33][17].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[33][17].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[33][17].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[33][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[33][17].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[33][18].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[33][18].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[33][18].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[33][18].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[33][18].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[33][18].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[33][18].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[33][18].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[33][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[33][18].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[33][19].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[33][19].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[33][19].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[33][19].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[33][19].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[33][19].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[33][19].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[33][19].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[33][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[33][19].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[33][20].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[33][20].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[33][20].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[33][20].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[33][20].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[33][20].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[33][20].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[33][20].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[33][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[33][20].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[33][21].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[33][21].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[33][21].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[33][21].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[33][21].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[33][21].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[33][21].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[33][21].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[33][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[33][21].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[33][22].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[33][22].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[33][22].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[33][22].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[33][22].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[33][22].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[33][22].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[33][22].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[33][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[33][22].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[33][23].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[33][23].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[33][23].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[33][23].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[33][23].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[33][23].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[33][23].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[33][23].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[33][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[33][23].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[33][24].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[33][24].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[33][24].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[33][24].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[33][24].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[33][24].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[33][24].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[33][24].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[33][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[33][24].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[33][25].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[33][25].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[33][25].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[33][25].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[33][25].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[33][25].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[33][25].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[33][25].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[33][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[33][25].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[33][26].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[33][26].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[33][26].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[33][26].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[33][26].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[33][26].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[33][26].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[33][26].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[33][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[33][26].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[33][27].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[33][27].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[33][27].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[33][27].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[33][27].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[33][27].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[33][27].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[33][27].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[33][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[33][27].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[33][28].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[33][28].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[33][28].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[33][28].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[33][28].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[33][28].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[33][28].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[33][28].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[33][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[33][28].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[33][29].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[33][29].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[33][29].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[33][29].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[33][29].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[33][29].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[33][29].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[33][29].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[33][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[33][29].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[33][30].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[33][30].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[33][30].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[33][30].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[33][30].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[33][30].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[33][30].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[33][30].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[33][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[33][30].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[33][31].dma__memc__write_valid      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[33][31].dma__memc__write_address    = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[33][31].dma__memc__write_data       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[33][31].dma__memc__read_valid       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[33][31].dma__memc__read_address     = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[33][31].dma__memc__read_pause       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[33][31].memc__dma__write_ready      = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[33][31].memc__dma__read_data        = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[33][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[33][31].memc__dma__read_ready       = pe_array_inst.pe_inst[33].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 34
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[34][0].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[34][0].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[34][0].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[34][0].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[34][0].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[34][0].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[34][0].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[34][0].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[34][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[34][0].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[34][1].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[34][1].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[34][1].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[34][1].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[34][1].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[34][1].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[34][1].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[34][1].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[34][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[34][1].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[34][2].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[34][2].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[34][2].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[34][2].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[34][2].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[34][2].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[34][2].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[34][2].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[34][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[34][2].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[34][3].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[34][3].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[34][3].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[34][3].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[34][3].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[34][3].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[34][3].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[34][3].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[34][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[34][3].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[34][4].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[34][4].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[34][4].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[34][4].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[34][4].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[34][4].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[34][4].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[34][4].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[34][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[34][4].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[34][5].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[34][5].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[34][5].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[34][5].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[34][5].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[34][5].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[34][5].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[34][5].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[34][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[34][5].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[34][6].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[34][6].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[34][6].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[34][6].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[34][6].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[34][6].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[34][6].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[34][6].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[34][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[34][6].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[34][7].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[34][7].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[34][7].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[34][7].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[34][7].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[34][7].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[34][7].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[34][7].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[34][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[34][7].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[34][8].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[34][8].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[34][8].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[34][8].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[34][8].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[34][8].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[34][8].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[34][8].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[34][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[34][8].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[34][9].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[34][9].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[34][9].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[34][9].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[34][9].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[34][9].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[34][9].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[34][9].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[34][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[34][9].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[34][10].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[34][10].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[34][10].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[34][10].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[34][10].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[34][10].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[34][10].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[34][10].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[34][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[34][10].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[34][11].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[34][11].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[34][11].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[34][11].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[34][11].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[34][11].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[34][11].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[34][11].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[34][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[34][11].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[34][12].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[34][12].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[34][12].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[34][12].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[34][12].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[34][12].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[34][12].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[34][12].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[34][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[34][12].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[34][13].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[34][13].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[34][13].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[34][13].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[34][13].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[34][13].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[34][13].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[34][13].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[34][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[34][13].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[34][14].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[34][14].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[34][14].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[34][14].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[34][14].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[34][14].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[34][14].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[34][14].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[34][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[34][14].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[34][15].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[34][15].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[34][15].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[34][15].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[34][15].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[34][15].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[34][15].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[34][15].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[34][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[34][15].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[34][16].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[34][16].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[34][16].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[34][16].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[34][16].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[34][16].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[34][16].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[34][16].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[34][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[34][16].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[34][17].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[34][17].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[34][17].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[34][17].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[34][17].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[34][17].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[34][17].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[34][17].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[34][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[34][17].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[34][18].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[34][18].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[34][18].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[34][18].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[34][18].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[34][18].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[34][18].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[34][18].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[34][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[34][18].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[34][19].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[34][19].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[34][19].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[34][19].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[34][19].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[34][19].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[34][19].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[34][19].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[34][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[34][19].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[34][20].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[34][20].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[34][20].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[34][20].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[34][20].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[34][20].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[34][20].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[34][20].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[34][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[34][20].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[34][21].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[34][21].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[34][21].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[34][21].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[34][21].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[34][21].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[34][21].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[34][21].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[34][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[34][21].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[34][22].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[34][22].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[34][22].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[34][22].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[34][22].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[34][22].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[34][22].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[34][22].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[34][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[34][22].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[34][23].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[34][23].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[34][23].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[34][23].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[34][23].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[34][23].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[34][23].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[34][23].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[34][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[34][23].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[34][24].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[34][24].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[34][24].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[34][24].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[34][24].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[34][24].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[34][24].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[34][24].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[34][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[34][24].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[34][25].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[34][25].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[34][25].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[34][25].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[34][25].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[34][25].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[34][25].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[34][25].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[34][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[34][25].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[34][26].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[34][26].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[34][26].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[34][26].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[34][26].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[34][26].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[34][26].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[34][26].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[34][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[34][26].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[34][27].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[34][27].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[34][27].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[34][27].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[34][27].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[34][27].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[34][27].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[34][27].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[34][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[34][27].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[34][28].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[34][28].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[34][28].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[34][28].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[34][28].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[34][28].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[34][28].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[34][28].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[34][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[34][28].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[34][29].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[34][29].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[34][29].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[34][29].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[34][29].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[34][29].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[34][29].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[34][29].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[34][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[34][29].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[34][30].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[34][30].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[34][30].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[34][30].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[34][30].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[34][30].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[34][30].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[34][30].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[34][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[34][30].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[34][31].dma__memc__write_valid      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[34][31].dma__memc__write_address    = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[34][31].dma__memc__write_data       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[34][31].dma__memc__read_valid       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[34][31].dma__memc__read_address     = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[34][31].dma__memc__read_pause       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[34][31].memc__dma__write_ready      = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[34][31].memc__dma__read_data        = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[34][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[34][31].memc__dma__read_ready       = pe_array_inst.pe_inst[34].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 35
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[35][0].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[35][0].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[35][0].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[35][0].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[35][0].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[35][0].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[35][0].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[35][0].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[35][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[35][0].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[35][1].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[35][1].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[35][1].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[35][1].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[35][1].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[35][1].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[35][1].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[35][1].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[35][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[35][1].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[35][2].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[35][2].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[35][2].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[35][2].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[35][2].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[35][2].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[35][2].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[35][2].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[35][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[35][2].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[35][3].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[35][3].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[35][3].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[35][3].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[35][3].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[35][3].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[35][3].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[35][3].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[35][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[35][3].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[35][4].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[35][4].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[35][4].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[35][4].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[35][4].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[35][4].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[35][4].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[35][4].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[35][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[35][4].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[35][5].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[35][5].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[35][5].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[35][5].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[35][5].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[35][5].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[35][5].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[35][5].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[35][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[35][5].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[35][6].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[35][6].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[35][6].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[35][6].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[35][6].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[35][6].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[35][6].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[35][6].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[35][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[35][6].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[35][7].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[35][7].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[35][7].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[35][7].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[35][7].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[35][7].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[35][7].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[35][7].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[35][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[35][7].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[35][8].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[35][8].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[35][8].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[35][8].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[35][8].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[35][8].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[35][8].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[35][8].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[35][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[35][8].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[35][9].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[35][9].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[35][9].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[35][9].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[35][9].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[35][9].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[35][9].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[35][9].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[35][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[35][9].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[35][10].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[35][10].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[35][10].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[35][10].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[35][10].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[35][10].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[35][10].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[35][10].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[35][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[35][10].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[35][11].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[35][11].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[35][11].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[35][11].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[35][11].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[35][11].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[35][11].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[35][11].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[35][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[35][11].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[35][12].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[35][12].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[35][12].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[35][12].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[35][12].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[35][12].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[35][12].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[35][12].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[35][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[35][12].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[35][13].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[35][13].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[35][13].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[35][13].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[35][13].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[35][13].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[35][13].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[35][13].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[35][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[35][13].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[35][14].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[35][14].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[35][14].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[35][14].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[35][14].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[35][14].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[35][14].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[35][14].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[35][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[35][14].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[35][15].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[35][15].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[35][15].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[35][15].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[35][15].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[35][15].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[35][15].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[35][15].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[35][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[35][15].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[35][16].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[35][16].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[35][16].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[35][16].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[35][16].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[35][16].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[35][16].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[35][16].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[35][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[35][16].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[35][17].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[35][17].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[35][17].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[35][17].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[35][17].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[35][17].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[35][17].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[35][17].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[35][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[35][17].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[35][18].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[35][18].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[35][18].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[35][18].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[35][18].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[35][18].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[35][18].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[35][18].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[35][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[35][18].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[35][19].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[35][19].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[35][19].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[35][19].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[35][19].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[35][19].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[35][19].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[35][19].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[35][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[35][19].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[35][20].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[35][20].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[35][20].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[35][20].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[35][20].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[35][20].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[35][20].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[35][20].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[35][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[35][20].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[35][21].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[35][21].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[35][21].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[35][21].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[35][21].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[35][21].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[35][21].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[35][21].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[35][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[35][21].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[35][22].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[35][22].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[35][22].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[35][22].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[35][22].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[35][22].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[35][22].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[35][22].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[35][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[35][22].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[35][23].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[35][23].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[35][23].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[35][23].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[35][23].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[35][23].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[35][23].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[35][23].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[35][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[35][23].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[35][24].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[35][24].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[35][24].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[35][24].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[35][24].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[35][24].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[35][24].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[35][24].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[35][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[35][24].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[35][25].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[35][25].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[35][25].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[35][25].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[35][25].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[35][25].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[35][25].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[35][25].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[35][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[35][25].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[35][26].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[35][26].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[35][26].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[35][26].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[35][26].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[35][26].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[35][26].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[35][26].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[35][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[35][26].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[35][27].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[35][27].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[35][27].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[35][27].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[35][27].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[35][27].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[35][27].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[35][27].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[35][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[35][27].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[35][28].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[35][28].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[35][28].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[35][28].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[35][28].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[35][28].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[35][28].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[35][28].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[35][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[35][28].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[35][29].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[35][29].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[35][29].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[35][29].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[35][29].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[35][29].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[35][29].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[35][29].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[35][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[35][29].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[35][30].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[35][30].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[35][30].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[35][30].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[35][30].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[35][30].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[35][30].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[35][30].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[35][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[35][30].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[35][31].dma__memc__write_valid      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[35][31].dma__memc__write_address    = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[35][31].dma__memc__write_data       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[35][31].dma__memc__read_valid       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[35][31].dma__memc__read_address     = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[35][31].dma__memc__read_pause       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[35][31].memc__dma__write_ready      = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[35][31].memc__dma__read_data        = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[35][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[35][31].memc__dma__read_ready       = pe_array_inst.pe_inst[35].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 36
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[36][0].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[36][0].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[36][0].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[36][0].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[36][0].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[36][0].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[36][0].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[36][0].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[36][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[36][0].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[36][1].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[36][1].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[36][1].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[36][1].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[36][1].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[36][1].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[36][1].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[36][1].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[36][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[36][1].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[36][2].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[36][2].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[36][2].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[36][2].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[36][2].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[36][2].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[36][2].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[36][2].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[36][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[36][2].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[36][3].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[36][3].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[36][3].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[36][3].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[36][3].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[36][3].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[36][3].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[36][3].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[36][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[36][3].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[36][4].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[36][4].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[36][4].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[36][4].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[36][4].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[36][4].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[36][4].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[36][4].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[36][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[36][4].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[36][5].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[36][5].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[36][5].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[36][5].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[36][5].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[36][5].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[36][5].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[36][5].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[36][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[36][5].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[36][6].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[36][6].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[36][6].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[36][6].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[36][6].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[36][6].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[36][6].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[36][6].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[36][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[36][6].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[36][7].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[36][7].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[36][7].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[36][7].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[36][7].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[36][7].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[36][7].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[36][7].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[36][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[36][7].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[36][8].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[36][8].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[36][8].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[36][8].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[36][8].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[36][8].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[36][8].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[36][8].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[36][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[36][8].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[36][9].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[36][9].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[36][9].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[36][9].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[36][9].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[36][9].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[36][9].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[36][9].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[36][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[36][9].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[36][10].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[36][10].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[36][10].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[36][10].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[36][10].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[36][10].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[36][10].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[36][10].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[36][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[36][10].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[36][11].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[36][11].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[36][11].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[36][11].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[36][11].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[36][11].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[36][11].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[36][11].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[36][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[36][11].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[36][12].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[36][12].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[36][12].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[36][12].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[36][12].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[36][12].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[36][12].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[36][12].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[36][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[36][12].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[36][13].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[36][13].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[36][13].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[36][13].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[36][13].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[36][13].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[36][13].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[36][13].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[36][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[36][13].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[36][14].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[36][14].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[36][14].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[36][14].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[36][14].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[36][14].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[36][14].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[36][14].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[36][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[36][14].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[36][15].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[36][15].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[36][15].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[36][15].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[36][15].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[36][15].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[36][15].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[36][15].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[36][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[36][15].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[36][16].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[36][16].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[36][16].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[36][16].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[36][16].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[36][16].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[36][16].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[36][16].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[36][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[36][16].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[36][17].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[36][17].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[36][17].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[36][17].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[36][17].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[36][17].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[36][17].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[36][17].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[36][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[36][17].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[36][18].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[36][18].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[36][18].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[36][18].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[36][18].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[36][18].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[36][18].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[36][18].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[36][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[36][18].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[36][19].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[36][19].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[36][19].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[36][19].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[36][19].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[36][19].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[36][19].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[36][19].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[36][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[36][19].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[36][20].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[36][20].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[36][20].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[36][20].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[36][20].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[36][20].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[36][20].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[36][20].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[36][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[36][20].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[36][21].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[36][21].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[36][21].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[36][21].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[36][21].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[36][21].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[36][21].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[36][21].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[36][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[36][21].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[36][22].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[36][22].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[36][22].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[36][22].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[36][22].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[36][22].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[36][22].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[36][22].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[36][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[36][22].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[36][23].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[36][23].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[36][23].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[36][23].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[36][23].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[36][23].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[36][23].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[36][23].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[36][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[36][23].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[36][24].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[36][24].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[36][24].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[36][24].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[36][24].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[36][24].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[36][24].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[36][24].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[36][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[36][24].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[36][25].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[36][25].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[36][25].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[36][25].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[36][25].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[36][25].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[36][25].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[36][25].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[36][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[36][25].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[36][26].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[36][26].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[36][26].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[36][26].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[36][26].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[36][26].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[36][26].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[36][26].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[36][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[36][26].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[36][27].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[36][27].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[36][27].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[36][27].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[36][27].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[36][27].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[36][27].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[36][27].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[36][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[36][27].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[36][28].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[36][28].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[36][28].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[36][28].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[36][28].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[36][28].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[36][28].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[36][28].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[36][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[36][28].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[36][29].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[36][29].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[36][29].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[36][29].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[36][29].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[36][29].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[36][29].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[36][29].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[36][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[36][29].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[36][30].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[36][30].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[36][30].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[36][30].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[36][30].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[36][30].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[36][30].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[36][30].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[36][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[36][30].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[36][31].dma__memc__write_valid      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[36][31].dma__memc__write_address    = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[36][31].dma__memc__write_data       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[36][31].dma__memc__read_valid       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[36][31].dma__memc__read_address     = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[36][31].dma__memc__read_pause       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[36][31].memc__dma__write_ready      = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[36][31].memc__dma__read_data        = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[36][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[36][31].memc__dma__read_ready       = pe_array_inst.pe_inst[36].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 37
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[37][0].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[37][0].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[37][0].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[37][0].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[37][0].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[37][0].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[37][0].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[37][0].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[37][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[37][0].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[37][1].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[37][1].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[37][1].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[37][1].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[37][1].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[37][1].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[37][1].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[37][1].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[37][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[37][1].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[37][2].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[37][2].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[37][2].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[37][2].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[37][2].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[37][2].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[37][2].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[37][2].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[37][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[37][2].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[37][3].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[37][3].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[37][3].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[37][3].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[37][3].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[37][3].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[37][3].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[37][3].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[37][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[37][3].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[37][4].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[37][4].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[37][4].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[37][4].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[37][4].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[37][4].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[37][4].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[37][4].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[37][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[37][4].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[37][5].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[37][5].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[37][5].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[37][5].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[37][5].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[37][5].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[37][5].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[37][5].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[37][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[37][5].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[37][6].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[37][6].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[37][6].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[37][6].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[37][6].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[37][6].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[37][6].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[37][6].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[37][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[37][6].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[37][7].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[37][7].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[37][7].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[37][7].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[37][7].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[37][7].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[37][7].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[37][7].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[37][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[37][7].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[37][8].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[37][8].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[37][8].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[37][8].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[37][8].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[37][8].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[37][8].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[37][8].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[37][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[37][8].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[37][9].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[37][9].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[37][9].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[37][9].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[37][9].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[37][9].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[37][9].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[37][9].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[37][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[37][9].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[37][10].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[37][10].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[37][10].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[37][10].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[37][10].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[37][10].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[37][10].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[37][10].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[37][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[37][10].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[37][11].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[37][11].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[37][11].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[37][11].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[37][11].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[37][11].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[37][11].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[37][11].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[37][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[37][11].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[37][12].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[37][12].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[37][12].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[37][12].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[37][12].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[37][12].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[37][12].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[37][12].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[37][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[37][12].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[37][13].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[37][13].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[37][13].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[37][13].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[37][13].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[37][13].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[37][13].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[37][13].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[37][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[37][13].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[37][14].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[37][14].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[37][14].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[37][14].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[37][14].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[37][14].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[37][14].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[37][14].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[37][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[37][14].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[37][15].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[37][15].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[37][15].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[37][15].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[37][15].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[37][15].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[37][15].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[37][15].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[37][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[37][15].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[37][16].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[37][16].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[37][16].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[37][16].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[37][16].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[37][16].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[37][16].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[37][16].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[37][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[37][16].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[37][17].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[37][17].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[37][17].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[37][17].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[37][17].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[37][17].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[37][17].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[37][17].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[37][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[37][17].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[37][18].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[37][18].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[37][18].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[37][18].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[37][18].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[37][18].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[37][18].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[37][18].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[37][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[37][18].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[37][19].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[37][19].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[37][19].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[37][19].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[37][19].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[37][19].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[37][19].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[37][19].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[37][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[37][19].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[37][20].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[37][20].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[37][20].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[37][20].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[37][20].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[37][20].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[37][20].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[37][20].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[37][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[37][20].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[37][21].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[37][21].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[37][21].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[37][21].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[37][21].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[37][21].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[37][21].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[37][21].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[37][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[37][21].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[37][22].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[37][22].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[37][22].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[37][22].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[37][22].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[37][22].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[37][22].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[37][22].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[37][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[37][22].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[37][23].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[37][23].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[37][23].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[37][23].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[37][23].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[37][23].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[37][23].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[37][23].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[37][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[37][23].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[37][24].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[37][24].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[37][24].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[37][24].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[37][24].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[37][24].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[37][24].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[37][24].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[37][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[37][24].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[37][25].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[37][25].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[37][25].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[37][25].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[37][25].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[37][25].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[37][25].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[37][25].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[37][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[37][25].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[37][26].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[37][26].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[37][26].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[37][26].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[37][26].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[37][26].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[37][26].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[37][26].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[37][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[37][26].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[37][27].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[37][27].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[37][27].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[37][27].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[37][27].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[37][27].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[37][27].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[37][27].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[37][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[37][27].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[37][28].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[37][28].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[37][28].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[37][28].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[37][28].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[37][28].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[37][28].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[37][28].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[37][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[37][28].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[37][29].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[37][29].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[37][29].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[37][29].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[37][29].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[37][29].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[37][29].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[37][29].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[37][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[37][29].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[37][30].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[37][30].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[37][30].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[37][30].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[37][30].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[37][30].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[37][30].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[37][30].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[37][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[37][30].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[37][31].dma__memc__write_valid      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[37][31].dma__memc__write_address    = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[37][31].dma__memc__write_data       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[37][31].dma__memc__read_valid       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[37][31].dma__memc__read_address     = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[37][31].dma__memc__read_pause       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[37][31].memc__dma__write_ready      = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[37][31].memc__dma__read_data        = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[37][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[37][31].memc__dma__read_ready       = pe_array_inst.pe_inst[37].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 38
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[38][0].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[38][0].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[38][0].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[38][0].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[38][0].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[38][0].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[38][0].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[38][0].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[38][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[38][0].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[38][1].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[38][1].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[38][1].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[38][1].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[38][1].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[38][1].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[38][1].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[38][1].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[38][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[38][1].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[38][2].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[38][2].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[38][2].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[38][2].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[38][2].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[38][2].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[38][2].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[38][2].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[38][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[38][2].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[38][3].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[38][3].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[38][3].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[38][3].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[38][3].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[38][3].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[38][3].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[38][3].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[38][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[38][3].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[38][4].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[38][4].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[38][4].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[38][4].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[38][4].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[38][4].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[38][4].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[38][4].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[38][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[38][4].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[38][5].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[38][5].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[38][5].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[38][5].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[38][5].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[38][5].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[38][5].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[38][5].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[38][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[38][5].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[38][6].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[38][6].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[38][6].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[38][6].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[38][6].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[38][6].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[38][6].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[38][6].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[38][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[38][6].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[38][7].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[38][7].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[38][7].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[38][7].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[38][7].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[38][7].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[38][7].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[38][7].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[38][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[38][7].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[38][8].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[38][8].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[38][8].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[38][8].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[38][8].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[38][8].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[38][8].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[38][8].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[38][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[38][8].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[38][9].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[38][9].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[38][9].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[38][9].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[38][9].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[38][9].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[38][9].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[38][9].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[38][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[38][9].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[38][10].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[38][10].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[38][10].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[38][10].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[38][10].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[38][10].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[38][10].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[38][10].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[38][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[38][10].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[38][11].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[38][11].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[38][11].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[38][11].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[38][11].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[38][11].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[38][11].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[38][11].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[38][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[38][11].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[38][12].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[38][12].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[38][12].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[38][12].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[38][12].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[38][12].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[38][12].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[38][12].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[38][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[38][12].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[38][13].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[38][13].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[38][13].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[38][13].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[38][13].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[38][13].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[38][13].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[38][13].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[38][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[38][13].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[38][14].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[38][14].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[38][14].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[38][14].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[38][14].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[38][14].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[38][14].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[38][14].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[38][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[38][14].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[38][15].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[38][15].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[38][15].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[38][15].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[38][15].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[38][15].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[38][15].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[38][15].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[38][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[38][15].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[38][16].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[38][16].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[38][16].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[38][16].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[38][16].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[38][16].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[38][16].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[38][16].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[38][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[38][16].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[38][17].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[38][17].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[38][17].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[38][17].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[38][17].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[38][17].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[38][17].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[38][17].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[38][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[38][17].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[38][18].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[38][18].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[38][18].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[38][18].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[38][18].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[38][18].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[38][18].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[38][18].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[38][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[38][18].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[38][19].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[38][19].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[38][19].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[38][19].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[38][19].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[38][19].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[38][19].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[38][19].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[38][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[38][19].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[38][20].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[38][20].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[38][20].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[38][20].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[38][20].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[38][20].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[38][20].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[38][20].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[38][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[38][20].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[38][21].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[38][21].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[38][21].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[38][21].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[38][21].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[38][21].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[38][21].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[38][21].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[38][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[38][21].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[38][22].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[38][22].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[38][22].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[38][22].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[38][22].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[38][22].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[38][22].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[38][22].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[38][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[38][22].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[38][23].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[38][23].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[38][23].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[38][23].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[38][23].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[38][23].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[38][23].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[38][23].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[38][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[38][23].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[38][24].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[38][24].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[38][24].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[38][24].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[38][24].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[38][24].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[38][24].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[38][24].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[38][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[38][24].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[38][25].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[38][25].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[38][25].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[38][25].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[38][25].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[38][25].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[38][25].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[38][25].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[38][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[38][25].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[38][26].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[38][26].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[38][26].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[38][26].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[38][26].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[38][26].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[38][26].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[38][26].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[38][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[38][26].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[38][27].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[38][27].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[38][27].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[38][27].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[38][27].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[38][27].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[38][27].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[38][27].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[38][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[38][27].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[38][28].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[38][28].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[38][28].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[38][28].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[38][28].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[38][28].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[38][28].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[38][28].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[38][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[38][28].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[38][29].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[38][29].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[38][29].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[38][29].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[38][29].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[38][29].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[38][29].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[38][29].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[38][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[38][29].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[38][30].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[38][30].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[38][30].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[38][30].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[38][30].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[38][30].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[38][30].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[38][30].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[38][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[38][30].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[38][31].dma__memc__write_valid      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[38][31].dma__memc__write_address    = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[38][31].dma__memc__write_data       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[38][31].dma__memc__read_valid       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[38][31].dma__memc__read_address     = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[38][31].dma__memc__read_pause       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[38][31].memc__dma__write_ready      = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[38][31].memc__dma__read_data        = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[38][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[38][31].memc__dma__read_ready       = pe_array_inst.pe_inst[38].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 39
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[39][0].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[39][0].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[39][0].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[39][0].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[39][0].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[39][0].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[39][0].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[39][0].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[39][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[39][0].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[39][1].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[39][1].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[39][1].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[39][1].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[39][1].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[39][1].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[39][1].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[39][1].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[39][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[39][1].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[39][2].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[39][2].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[39][2].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[39][2].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[39][2].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[39][2].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[39][2].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[39][2].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[39][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[39][2].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[39][3].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[39][3].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[39][3].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[39][3].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[39][3].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[39][3].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[39][3].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[39][3].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[39][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[39][3].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[39][4].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[39][4].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[39][4].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[39][4].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[39][4].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[39][4].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[39][4].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[39][4].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[39][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[39][4].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[39][5].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[39][5].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[39][5].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[39][5].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[39][5].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[39][5].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[39][5].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[39][5].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[39][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[39][5].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[39][6].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[39][6].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[39][6].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[39][6].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[39][6].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[39][6].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[39][6].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[39][6].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[39][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[39][6].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[39][7].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[39][7].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[39][7].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[39][7].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[39][7].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[39][7].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[39][7].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[39][7].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[39][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[39][7].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[39][8].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[39][8].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[39][8].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[39][8].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[39][8].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[39][8].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[39][8].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[39][8].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[39][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[39][8].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[39][9].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[39][9].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[39][9].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[39][9].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[39][9].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[39][9].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[39][9].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[39][9].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[39][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[39][9].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[39][10].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[39][10].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[39][10].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[39][10].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[39][10].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[39][10].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[39][10].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[39][10].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[39][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[39][10].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[39][11].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[39][11].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[39][11].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[39][11].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[39][11].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[39][11].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[39][11].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[39][11].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[39][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[39][11].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[39][12].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[39][12].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[39][12].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[39][12].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[39][12].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[39][12].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[39][12].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[39][12].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[39][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[39][12].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[39][13].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[39][13].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[39][13].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[39][13].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[39][13].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[39][13].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[39][13].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[39][13].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[39][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[39][13].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[39][14].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[39][14].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[39][14].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[39][14].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[39][14].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[39][14].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[39][14].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[39][14].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[39][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[39][14].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[39][15].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[39][15].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[39][15].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[39][15].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[39][15].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[39][15].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[39][15].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[39][15].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[39][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[39][15].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[39][16].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[39][16].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[39][16].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[39][16].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[39][16].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[39][16].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[39][16].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[39][16].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[39][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[39][16].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[39][17].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[39][17].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[39][17].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[39][17].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[39][17].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[39][17].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[39][17].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[39][17].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[39][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[39][17].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[39][18].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[39][18].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[39][18].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[39][18].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[39][18].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[39][18].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[39][18].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[39][18].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[39][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[39][18].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[39][19].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[39][19].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[39][19].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[39][19].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[39][19].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[39][19].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[39][19].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[39][19].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[39][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[39][19].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[39][20].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[39][20].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[39][20].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[39][20].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[39][20].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[39][20].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[39][20].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[39][20].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[39][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[39][20].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[39][21].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[39][21].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[39][21].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[39][21].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[39][21].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[39][21].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[39][21].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[39][21].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[39][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[39][21].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[39][22].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[39][22].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[39][22].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[39][22].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[39][22].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[39][22].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[39][22].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[39][22].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[39][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[39][22].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[39][23].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[39][23].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[39][23].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[39][23].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[39][23].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[39][23].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[39][23].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[39][23].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[39][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[39][23].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[39][24].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[39][24].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[39][24].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[39][24].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[39][24].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[39][24].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[39][24].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[39][24].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[39][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[39][24].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[39][25].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[39][25].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[39][25].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[39][25].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[39][25].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[39][25].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[39][25].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[39][25].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[39][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[39][25].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[39][26].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[39][26].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[39][26].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[39][26].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[39][26].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[39][26].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[39][26].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[39][26].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[39][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[39][26].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[39][27].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[39][27].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[39][27].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[39][27].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[39][27].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[39][27].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[39][27].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[39][27].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[39][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[39][27].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[39][28].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[39][28].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[39][28].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[39][28].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[39][28].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[39][28].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[39][28].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[39][28].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[39][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[39][28].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[39][29].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[39][29].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[39][29].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[39][29].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[39][29].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[39][29].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[39][29].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[39][29].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[39][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[39][29].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[39][30].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[39][30].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[39][30].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[39][30].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[39][30].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[39][30].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[39][30].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[39][30].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[39][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[39][30].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[39][31].dma__memc__write_valid      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[39][31].dma__memc__write_address    = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[39][31].dma__memc__write_data       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[39][31].dma__memc__read_valid       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[39][31].dma__memc__read_address     = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[39][31].dma__memc__read_pause       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[39][31].memc__dma__write_ready      = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[39][31].memc__dma__read_data        = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[39][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[39][31].memc__dma__read_ready       = pe_array_inst.pe_inst[39].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 40
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[40][0].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[40][0].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[40][0].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[40][0].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[40][0].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[40][0].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[40][0].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[40][0].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[40][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[40][0].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[40][1].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[40][1].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[40][1].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[40][1].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[40][1].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[40][1].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[40][1].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[40][1].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[40][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[40][1].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[40][2].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[40][2].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[40][2].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[40][2].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[40][2].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[40][2].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[40][2].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[40][2].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[40][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[40][2].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[40][3].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[40][3].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[40][3].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[40][3].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[40][3].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[40][3].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[40][3].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[40][3].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[40][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[40][3].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[40][4].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[40][4].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[40][4].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[40][4].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[40][4].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[40][4].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[40][4].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[40][4].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[40][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[40][4].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[40][5].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[40][5].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[40][5].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[40][5].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[40][5].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[40][5].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[40][5].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[40][5].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[40][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[40][5].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[40][6].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[40][6].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[40][6].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[40][6].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[40][6].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[40][6].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[40][6].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[40][6].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[40][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[40][6].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[40][7].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[40][7].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[40][7].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[40][7].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[40][7].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[40][7].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[40][7].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[40][7].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[40][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[40][7].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[40][8].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[40][8].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[40][8].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[40][8].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[40][8].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[40][8].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[40][8].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[40][8].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[40][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[40][8].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[40][9].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[40][9].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[40][9].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[40][9].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[40][9].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[40][9].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[40][9].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[40][9].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[40][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[40][9].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[40][10].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[40][10].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[40][10].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[40][10].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[40][10].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[40][10].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[40][10].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[40][10].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[40][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[40][10].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[40][11].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[40][11].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[40][11].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[40][11].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[40][11].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[40][11].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[40][11].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[40][11].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[40][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[40][11].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[40][12].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[40][12].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[40][12].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[40][12].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[40][12].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[40][12].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[40][12].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[40][12].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[40][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[40][12].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[40][13].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[40][13].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[40][13].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[40][13].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[40][13].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[40][13].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[40][13].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[40][13].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[40][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[40][13].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[40][14].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[40][14].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[40][14].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[40][14].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[40][14].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[40][14].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[40][14].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[40][14].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[40][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[40][14].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[40][15].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[40][15].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[40][15].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[40][15].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[40][15].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[40][15].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[40][15].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[40][15].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[40][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[40][15].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[40][16].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[40][16].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[40][16].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[40][16].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[40][16].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[40][16].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[40][16].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[40][16].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[40][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[40][16].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[40][17].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[40][17].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[40][17].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[40][17].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[40][17].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[40][17].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[40][17].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[40][17].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[40][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[40][17].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[40][18].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[40][18].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[40][18].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[40][18].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[40][18].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[40][18].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[40][18].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[40][18].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[40][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[40][18].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[40][19].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[40][19].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[40][19].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[40][19].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[40][19].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[40][19].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[40][19].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[40][19].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[40][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[40][19].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[40][20].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[40][20].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[40][20].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[40][20].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[40][20].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[40][20].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[40][20].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[40][20].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[40][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[40][20].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[40][21].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[40][21].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[40][21].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[40][21].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[40][21].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[40][21].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[40][21].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[40][21].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[40][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[40][21].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[40][22].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[40][22].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[40][22].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[40][22].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[40][22].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[40][22].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[40][22].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[40][22].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[40][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[40][22].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[40][23].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[40][23].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[40][23].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[40][23].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[40][23].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[40][23].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[40][23].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[40][23].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[40][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[40][23].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[40][24].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[40][24].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[40][24].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[40][24].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[40][24].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[40][24].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[40][24].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[40][24].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[40][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[40][24].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[40][25].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[40][25].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[40][25].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[40][25].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[40][25].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[40][25].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[40][25].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[40][25].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[40][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[40][25].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[40][26].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[40][26].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[40][26].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[40][26].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[40][26].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[40][26].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[40][26].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[40][26].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[40][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[40][26].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[40][27].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[40][27].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[40][27].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[40][27].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[40][27].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[40][27].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[40][27].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[40][27].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[40][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[40][27].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[40][28].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[40][28].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[40][28].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[40][28].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[40][28].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[40][28].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[40][28].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[40][28].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[40][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[40][28].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[40][29].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[40][29].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[40][29].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[40][29].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[40][29].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[40][29].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[40][29].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[40][29].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[40][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[40][29].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[40][30].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[40][30].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[40][30].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[40][30].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[40][30].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[40][30].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[40][30].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[40][30].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[40][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[40][30].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[40][31].dma__memc__write_valid      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[40][31].dma__memc__write_address    = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[40][31].dma__memc__write_data       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[40][31].dma__memc__read_valid       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[40][31].dma__memc__read_address     = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[40][31].dma__memc__read_pause       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[40][31].memc__dma__write_ready      = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[40][31].memc__dma__read_data        = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[40][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[40][31].memc__dma__read_ready       = pe_array_inst.pe_inst[40].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 41
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[41][0].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[41][0].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[41][0].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[41][0].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[41][0].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[41][0].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[41][0].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[41][0].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[41][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[41][0].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[41][1].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[41][1].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[41][1].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[41][1].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[41][1].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[41][1].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[41][1].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[41][1].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[41][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[41][1].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[41][2].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[41][2].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[41][2].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[41][2].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[41][2].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[41][2].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[41][2].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[41][2].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[41][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[41][2].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[41][3].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[41][3].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[41][3].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[41][3].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[41][3].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[41][3].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[41][3].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[41][3].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[41][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[41][3].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[41][4].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[41][4].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[41][4].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[41][4].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[41][4].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[41][4].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[41][4].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[41][4].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[41][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[41][4].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[41][5].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[41][5].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[41][5].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[41][5].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[41][5].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[41][5].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[41][5].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[41][5].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[41][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[41][5].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[41][6].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[41][6].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[41][6].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[41][6].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[41][6].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[41][6].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[41][6].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[41][6].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[41][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[41][6].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[41][7].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[41][7].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[41][7].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[41][7].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[41][7].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[41][7].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[41][7].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[41][7].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[41][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[41][7].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[41][8].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[41][8].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[41][8].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[41][8].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[41][8].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[41][8].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[41][8].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[41][8].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[41][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[41][8].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[41][9].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[41][9].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[41][9].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[41][9].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[41][9].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[41][9].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[41][9].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[41][9].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[41][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[41][9].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[41][10].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[41][10].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[41][10].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[41][10].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[41][10].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[41][10].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[41][10].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[41][10].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[41][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[41][10].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[41][11].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[41][11].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[41][11].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[41][11].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[41][11].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[41][11].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[41][11].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[41][11].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[41][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[41][11].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[41][12].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[41][12].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[41][12].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[41][12].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[41][12].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[41][12].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[41][12].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[41][12].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[41][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[41][12].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[41][13].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[41][13].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[41][13].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[41][13].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[41][13].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[41][13].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[41][13].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[41][13].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[41][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[41][13].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[41][14].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[41][14].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[41][14].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[41][14].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[41][14].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[41][14].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[41][14].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[41][14].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[41][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[41][14].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[41][15].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[41][15].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[41][15].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[41][15].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[41][15].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[41][15].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[41][15].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[41][15].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[41][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[41][15].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[41][16].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[41][16].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[41][16].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[41][16].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[41][16].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[41][16].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[41][16].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[41][16].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[41][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[41][16].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[41][17].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[41][17].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[41][17].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[41][17].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[41][17].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[41][17].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[41][17].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[41][17].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[41][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[41][17].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[41][18].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[41][18].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[41][18].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[41][18].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[41][18].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[41][18].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[41][18].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[41][18].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[41][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[41][18].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[41][19].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[41][19].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[41][19].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[41][19].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[41][19].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[41][19].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[41][19].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[41][19].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[41][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[41][19].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[41][20].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[41][20].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[41][20].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[41][20].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[41][20].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[41][20].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[41][20].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[41][20].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[41][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[41][20].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[41][21].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[41][21].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[41][21].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[41][21].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[41][21].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[41][21].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[41][21].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[41][21].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[41][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[41][21].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[41][22].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[41][22].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[41][22].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[41][22].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[41][22].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[41][22].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[41][22].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[41][22].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[41][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[41][22].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[41][23].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[41][23].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[41][23].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[41][23].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[41][23].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[41][23].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[41][23].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[41][23].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[41][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[41][23].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[41][24].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[41][24].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[41][24].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[41][24].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[41][24].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[41][24].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[41][24].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[41][24].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[41][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[41][24].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[41][25].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[41][25].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[41][25].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[41][25].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[41][25].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[41][25].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[41][25].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[41][25].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[41][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[41][25].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[41][26].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[41][26].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[41][26].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[41][26].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[41][26].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[41][26].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[41][26].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[41][26].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[41][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[41][26].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[41][27].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[41][27].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[41][27].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[41][27].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[41][27].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[41][27].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[41][27].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[41][27].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[41][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[41][27].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[41][28].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[41][28].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[41][28].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[41][28].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[41][28].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[41][28].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[41][28].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[41][28].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[41][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[41][28].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[41][29].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[41][29].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[41][29].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[41][29].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[41][29].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[41][29].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[41][29].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[41][29].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[41][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[41][29].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[41][30].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[41][30].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[41][30].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[41][30].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[41][30].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[41][30].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[41][30].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[41][30].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[41][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[41][30].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[41][31].dma__memc__write_valid      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[41][31].dma__memc__write_address    = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[41][31].dma__memc__write_data       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[41][31].dma__memc__read_valid       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[41][31].dma__memc__read_address     = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[41][31].dma__memc__read_pause       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[41][31].memc__dma__write_ready      = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[41][31].memc__dma__read_data        = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[41][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[41][31].memc__dma__read_ready       = pe_array_inst.pe_inst[41].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 42
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[42][0].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[42][0].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[42][0].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[42][0].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[42][0].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[42][0].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[42][0].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[42][0].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[42][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[42][0].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[42][1].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[42][1].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[42][1].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[42][1].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[42][1].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[42][1].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[42][1].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[42][1].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[42][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[42][1].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[42][2].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[42][2].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[42][2].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[42][2].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[42][2].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[42][2].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[42][2].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[42][2].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[42][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[42][2].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[42][3].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[42][3].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[42][3].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[42][3].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[42][3].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[42][3].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[42][3].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[42][3].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[42][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[42][3].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[42][4].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[42][4].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[42][4].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[42][4].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[42][4].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[42][4].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[42][4].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[42][4].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[42][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[42][4].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[42][5].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[42][5].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[42][5].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[42][5].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[42][5].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[42][5].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[42][5].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[42][5].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[42][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[42][5].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[42][6].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[42][6].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[42][6].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[42][6].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[42][6].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[42][6].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[42][6].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[42][6].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[42][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[42][6].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[42][7].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[42][7].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[42][7].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[42][7].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[42][7].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[42][7].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[42][7].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[42][7].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[42][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[42][7].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[42][8].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[42][8].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[42][8].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[42][8].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[42][8].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[42][8].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[42][8].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[42][8].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[42][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[42][8].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[42][9].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[42][9].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[42][9].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[42][9].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[42][9].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[42][9].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[42][9].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[42][9].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[42][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[42][9].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[42][10].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[42][10].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[42][10].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[42][10].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[42][10].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[42][10].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[42][10].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[42][10].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[42][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[42][10].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[42][11].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[42][11].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[42][11].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[42][11].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[42][11].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[42][11].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[42][11].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[42][11].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[42][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[42][11].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[42][12].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[42][12].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[42][12].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[42][12].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[42][12].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[42][12].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[42][12].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[42][12].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[42][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[42][12].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[42][13].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[42][13].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[42][13].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[42][13].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[42][13].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[42][13].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[42][13].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[42][13].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[42][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[42][13].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[42][14].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[42][14].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[42][14].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[42][14].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[42][14].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[42][14].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[42][14].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[42][14].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[42][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[42][14].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[42][15].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[42][15].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[42][15].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[42][15].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[42][15].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[42][15].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[42][15].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[42][15].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[42][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[42][15].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[42][16].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[42][16].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[42][16].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[42][16].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[42][16].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[42][16].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[42][16].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[42][16].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[42][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[42][16].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[42][17].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[42][17].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[42][17].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[42][17].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[42][17].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[42][17].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[42][17].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[42][17].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[42][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[42][17].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[42][18].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[42][18].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[42][18].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[42][18].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[42][18].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[42][18].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[42][18].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[42][18].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[42][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[42][18].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[42][19].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[42][19].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[42][19].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[42][19].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[42][19].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[42][19].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[42][19].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[42][19].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[42][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[42][19].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[42][20].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[42][20].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[42][20].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[42][20].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[42][20].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[42][20].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[42][20].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[42][20].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[42][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[42][20].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[42][21].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[42][21].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[42][21].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[42][21].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[42][21].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[42][21].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[42][21].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[42][21].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[42][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[42][21].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[42][22].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[42][22].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[42][22].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[42][22].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[42][22].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[42][22].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[42][22].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[42][22].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[42][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[42][22].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[42][23].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[42][23].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[42][23].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[42][23].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[42][23].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[42][23].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[42][23].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[42][23].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[42][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[42][23].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[42][24].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[42][24].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[42][24].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[42][24].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[42][24].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[42][24].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[42][24].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[42][24].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[42][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[42][24].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[42][25].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[42][25].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[42][25].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[42][25].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[42][25].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[42][25].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[42][25].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[42][25].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[42][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[42][25].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[42][26].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[42][26].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[42][26].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[42][26].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[42][26].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[42][26].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[42][26].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[42][26].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[42][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[42][26].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[42][27].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[42][27].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[42][27].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[42][27].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[42][27].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[42][27].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[42][27].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[42][27].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[42][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[42][27].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[42][28].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[42][28].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[42][28].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[42][28].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[42][28].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[42][28].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[42][28].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[42][28].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[42][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[42][28].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[42][29].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[42][29].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[42][29].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[42][29].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[42][29].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[42][29].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[42][29].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[42][29].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[42][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[42][29].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[42][30].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[42][30].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[42][30].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[42][30].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[42][30].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[42][30].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[42][30].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[42][30].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[42][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[42][30].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[42][31].dma__memc__write_valid      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[42][31].dma__memc__write_address    = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[42][31].dma__memc__write_data       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[42][31].dma__memc__read_valid       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[42][31].dma__memc__read_address     = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[42][31].dma__memc__read_pause       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[42][31].memc__dma__write_ready      = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[42][31].memc__dma__read_data        = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[42][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[42][31].memc__dma__read_ready       = pe_array_inst.pe_inst[42].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 43
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[43][0].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[43][0].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[43][0].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[43][0].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[43][0].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[43][0].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[43][0].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[43][0].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[43][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[43][0].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[43][1].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[43][1].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[43][1].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[43][1].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[43][1].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[43][1].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[43][1].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[43][1].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[43][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[43][1].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[43][2].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[43][2].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[43][2].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[43][2].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[43][2].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[43][2].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[43][2].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[43][2].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[43][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[43][2].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[43][3].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[43][3].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[43][3].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[43][3].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[43][3].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[43][3].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[43][3].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[43][3].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[43][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[43][3].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[43][4].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[43][4].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[43][4].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[43][4].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[43][4].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[43][4].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[43][4].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[43][4].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[43][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[43][4].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[43][5].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[43][5].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[43][5].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[43][5].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[43][5].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[43][5].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[43][5].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[43][5].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[43][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[43][5].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[43][6].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[43][6].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[43][6].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[43][6].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[43][6].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[43][6].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[43][6].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[43][6].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[43][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[43][6].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[43][7].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[43][7].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[43][7].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[43][7].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[43][7].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[43][7].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[43][7].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[43][7].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[43][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[43][7].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[43][8].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[43][8].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[43][8].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[43][8].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[43][8].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[43][8].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[43][8].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[43][8].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[43][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[43][8].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[43][9].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[43][9].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[43][9].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[43][9].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[43][9].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[43][9].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[43][9].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[43][9].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[43][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[43][9].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[43][10].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[43][10].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[43][10].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[43][10].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[43][10].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[43][10].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[43][10].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[43][10].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[43][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[43][10].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[43][11].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[43][11].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[43][11].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[43][11].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[43][11].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[43][11].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[43][11].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[43][11].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[43][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[43][11].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[43][12].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[43][12].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[43][12].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[43][12].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[43][12].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[43][12].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[43][12].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[43][12].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[43][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[43][12].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[43][13].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[43][13].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[43][13].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[43][13].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[43][13].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[43][13].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[43][13].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[43][13].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[43][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[43][13].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[43][14].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[43][14].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[43][14].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[43][14].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[43][14].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[43][14].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[43][14].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[43][14].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[43][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[43][14].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[43][15].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[43][15].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[43][15].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[43][15].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[43][15].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[43][15].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[43][15].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[43][15].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[43][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[43][15].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[43][16].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[43][16].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[43][16].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[43][16].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[43][16].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[43][16].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[43][16].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[43][16].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[43][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[43][16].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[43][17].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[43][17].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[43][17].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[43][17].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[43][17].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[43][17].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[43][17].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[43][17].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[43][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[43][17].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[43][18].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[43][18].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[43][18].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[43][18].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[43][18].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[43][18].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[43][18].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[43][18].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[43][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[43][18].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[43][19].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[43][19].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[43][19].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[43][19].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[43][19].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[43][19].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[43][19].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[43][19].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[43][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[43][19].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[43][20].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[43][20].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[43][20].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[43][20].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[43][20].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[43][20].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[43][20].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[43][20].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[43][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[43][20].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[43][21].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[43][21].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[43][21].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[43][21].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[43][21].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[43][21].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[43][21].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[43][21].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[43][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[43][21].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[43][22].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[43][22].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[43][22].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[43][22].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[43][22].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[43][22].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[43][22].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[43][22].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[43][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[43][22].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[43][23].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[43][23].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[43][23].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[43][23].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[43][23].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[43][23].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[43][23].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[43][23].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[43][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[43][23].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[43][24].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[43][24].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[43][24].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[43][24].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[43][24].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[43][24].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[43][24].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[43][24].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[43][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[43][24].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[43][25].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[43][25].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[43][25].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[43][25].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[43][25].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[43][25].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[43][25].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[43][25].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[43][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[43][25].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[43][26].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[43][26].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[43][26].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[43][26].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[43][26].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[43][26].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[43][26].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[43][26].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[43][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[43][26].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[43][27].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[43][27].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[43][27].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[43][27].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[43][27].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[43][27].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[43][27].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[43][27].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[43][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[43][27].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[43][28].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[43][28].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[43][28].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[43][28].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[43][28].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[43][28].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[43][28].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[43][28].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[43][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[43][28].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[43][29].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[43][29].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[43][29].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[43][29].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[43][29].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[43][29].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[43][29].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[43][29].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[43][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[43][29].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[43][30].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[43][30].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[43][30].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[43][30].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[43][30].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[43][30].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[43][30].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[43][30].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[43][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[43][30].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[43][31].dma__memc__write_valid      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[43][31].dma__memc__write_address    = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[43][31].dma__memc__write_data       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[43][31].dma__memc__read_valid       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[43][31].dma__memc__read_address     = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[43][31].dma__memc__read_pause       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[43][31].memc__dma__write_ready      = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[43][31].memc__dma__read_data        = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[43][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[43][31].memc__dma__read_ready       = pe_array_inst.pe_inst[43].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 44
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[44][0].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[44][0].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[44][0].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[44][0].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[44][0].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[44][0].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[44][0].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[44][0].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[44][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[44][0].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[44][1].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[44][1].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[44][1].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[44][1].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[44][1].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[44][1].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[44][1].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[44][1].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[44][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[44][1].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[44][2].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[44][2].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[44][2].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[44][2].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[44][2].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[44][2].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[44][2].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[44][2].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[44][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[44][2].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[44][3].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[44][3].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[44][3].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[44][3].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[44][3].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[44][3].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[44][3].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[44][3].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[44][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[44][3].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[44][4].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[44][4].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[44][4].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[44][4].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[44][4].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[44][4].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[44][4].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[44][4].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[44][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[44][4].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[44][5].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[44][5].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[44][5].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[44][5].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[44][5].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[44][5].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[44][5].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[44][5].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[44][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[44][5].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[44][6].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[44][6].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[44][6].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[44][6].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[44][6].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[44][6].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[44][6].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[44][6].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[44][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[44][6].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[44][7].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[44][7].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[44][7].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[44][7].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[44][7].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[44][7].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[44][7].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[44][7].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[44][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[44][7].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[44][8].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[44][8].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[44][8].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[44][8].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[44][8].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[44][8].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[44][8].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[44][8].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[44][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[44][8].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[44][9].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[44][9].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[44][9].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[44][9].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[44][9].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[44][9].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[44][9].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[44][9].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[44][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[44][9].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[44][10].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[44][10].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[44][10].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[44][10].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[44][10].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[44][10].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[44][10].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[44][10].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[44][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[44][10].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[44][11].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[44][11].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[44][11].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[44][11].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[44][11].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[44][11].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[44][11].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[44][11].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[44][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[44][11].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[44][12].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[44][12].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[44][12].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[44][12].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[44][12].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[44][12].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[44][12].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[44][12].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[44][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[44][12].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[44][13].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[44][13].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[44][13].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[44][13].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[44][13].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[44][13].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[44][13].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[44][13].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[44][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[44][13].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[44][14].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[44][14].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[44][14].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[44][14].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[44][14].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[44][14].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[44][14].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[44][14].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[44][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[44][14].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[44][15].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[44][15].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[44][15].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[44][15].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[44][15].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[44][15].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[44][15].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[44][15].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[44][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[44][15].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[44][16].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[44][16].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[44][16].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[44][16].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[44][16].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[44][16].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[44][16].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[44][16].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[44][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[44][16].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[44][17].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[44][17].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[44][17].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[44][17].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[44][17].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[44][17].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[44][17].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[44][17].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[44][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[44][17].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[44][18].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[44][18].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[44][18].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[44][18].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[44][18].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[44][18].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[44][18].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[44][18].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[44][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[44][18].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[44][19].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[44][19].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[44][19].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[44][19].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[44][19].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[44][19].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[44][19].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[44][19].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[44][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[44][19].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[44][20].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[44][20].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[44][20].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[44][20].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[44][20].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[44][20].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[44][20].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[44][20].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[44][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[44][20].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[44][21].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[44][21].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[44][21].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[44][21].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[44][21].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[44][21].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[44][21].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[44][21].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[44][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[44][21].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[44][22].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[44][22].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[44][22].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[44][22].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[44][22].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[44][22].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[44][22].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[44][22].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[44][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[44][22].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[44][23].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[44][23].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[44][23].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[44][23].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[44][23].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[44][23].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[44][23].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[44][23].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[44][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[44][23].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[44][24].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[44][24].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[44][24].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[44][24].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[44][24].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[44][24].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[44][24].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[44][24].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[44][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[44][24].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[44][25].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[44][25].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[44][25].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[44][25].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[44][25].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[44][25].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[44][25].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[44][25].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[44][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[44][25].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[44][26].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[44][26].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[44][26].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[44][26].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[44][26].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[44][26].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[44][26].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[44][26].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[44][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[44][26].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[44][27].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[44][27].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[44][27].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[44][27].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[44][27].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[44][27].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[44][27].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[44][27].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[44][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[44][27].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[44][28].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[44][28].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[44][28].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[44][28].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[44][28].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[44][28].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[44][28].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[44][28].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[44][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[44][28].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[44][29].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[44][29].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[44][29].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[44][29].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[44][29].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[44][29].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[44][29].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[44][29].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[44][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[44][29].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[44][30].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[44][30].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[44][30].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[44][30].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[44][30].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[44][30].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[44][30].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[44][30].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[44][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[44][30].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[44][31].dma__memc__write_valid      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[44][31].dma__memc__write_address    = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[44][31].dma__memc__write_data       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[44][31].dma__memc__read_valid       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[44][31].dma__memc__read_address     = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[44][31].dma__memc__read_pause       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[44][31].memc__dma__write_ready      = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[44][31].memc__dma__read_data        = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[44][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[44][31].memc__dma__read_ready       = pe_array_inst.pe_inst[44].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 45
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[45][0].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[45][0].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[45][0].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[45][0].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[45][0].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[45][0].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[45][0].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[45][0].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[45][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[45][0].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[45][1].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[45][1].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[45][1].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[45][1].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[45][1].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[45][1].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[45][1].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[45][1].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[45][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[45][1].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[45][2].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[45][2].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[45][2].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[45][2].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[45][2].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[45][2].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[45][2].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[45][2].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[45][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[45][2].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[45][3].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[45][3].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[45][3].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[45][3].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[45][3].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[45][3].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[45][3].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[45][3].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[45][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[45][3].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[45][4].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[45][4].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[45][4].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[45][4].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[45][4].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[45][4].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[45][4].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[45][4].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[45][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[45][4].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[45][5].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[45][5].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[45][5].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[45][5].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[45][5].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[45][5].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[45][5].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[45][5].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[45][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[45][5].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[45][6].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[45][6].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[45][6].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[45][6].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[45][6].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[45][6].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[45][6].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[45][6].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[45][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[45][6].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[45][7].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[45][7].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[45][7].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[45][7].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[45][7].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[45][7].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[45][7].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[45][7].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[45][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[45][7].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[45][8].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[45][8].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[45][8].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[45][8].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[45][8].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[45][8].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[45][8].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[45][8].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[45][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[45][8].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[45][9].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[45][9].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[45][9].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[45][9].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[45][9].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[45][9].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[45][9].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[45][9].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[45][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[45][9].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[45][10].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[45][10].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[45][10].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[45][10].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[45][10].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[45][10].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[45][10].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[45][10].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[45][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[45][10].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[45][11].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[45][11].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[45][11].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[45][11].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[45][11].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[45][11].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[45][11].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[45][11].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[45][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[45][11].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[45][12].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[45][12].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[45][12].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[45][12].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[45][12].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[45][12].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[45][12].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[45][12].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[45][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[45][12].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[45][13].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[45][13].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[45][13].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[45][13].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[45][13].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[45][13].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[45][13].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[45][13].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[45][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[45][13].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[45][14].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[45][14].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[45][14].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[45][14].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[45][14].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[45][14].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[45][14].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[45][14].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[45][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[45][14].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[45][15].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[45][15].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[45][15].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[45][15].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[45][15].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[45][15].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[45][15].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[45][15].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[45][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[45][15].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[45][16].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[45][16].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[45][16].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[45][16].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[45][16].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[45][16].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[45][16].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[45][16].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[45][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[45][16].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[45][17].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[45][17].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[45][17].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[45][17].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[45][17].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[45][17].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[45][17].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[45][17].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[45][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[45][17].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[45][18].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[45][18].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[45][18].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[45][18].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[45][18].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[45][18].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[45][18].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[45][18].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[45][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[45][18].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[45][19].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[45][19].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[45][19].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[45][19].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[45][19].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[45][19].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[45][19].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[45][19].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[45][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[45][19].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[45][20].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[45][20].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[45][20].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[45][20].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[45][20].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[45][20].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[45][20].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[45][20].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[45][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[45][20].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[45][21].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[45][21].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[45][21].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[45][21].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[45][21].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[45][21].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[45][21].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[45][21].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[45][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[45][21].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[45][22].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[45][22].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[45][22].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[45][22].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[45][22].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[45][22].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[45][22].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[45][22].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[45][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[45][22].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[45][23].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[45][23].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[45][23].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[45][23].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[45][23].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[45][23].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[45][23].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[45][23].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[45][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[45][23].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[45][24].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[45][24].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[45][24].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[45][24].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[45][24].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[45][24].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[45][24].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[45][24].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[45][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[45][24].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[45][25].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[45][25].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[45][25].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[45][25].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[45][25].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[45][25].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[45][25].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[45][25].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[45][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[45][25].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[45][26].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[45][26].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[45][26].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[45][26].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[45][26].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[45][26].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[45][26].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[45][26].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[45][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[45][26].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[45][27].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[45][27].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[45][27].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[45][27].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[45][27].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[45][27].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[45][27].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[45][27].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[45][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[45][27].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[45][28].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[45][28].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[45][28].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[45][28].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[45][28].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[45][28].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[45][28].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[45][28].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[45][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[45][28].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[45][29].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[45][29].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[45][29].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[45][29].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[45][29].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[45][29].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[45][29].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[45][29].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[45][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[45][29].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[45][30].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[45][30].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[45][30].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[45][30].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[45][30].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[45][30].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[45][30].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[45][30].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[45][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[45][30].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[45][31].dma__memc__write_valid      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[45][31].dma__memc__write_address    = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[45][31].dma__memc__write_data       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[45][31].dma__memc__read_valid       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[45][31].dma__memc__read_address     = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[45][31].dma__memc__read_pause       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[45][31].memc__dma__write_ready      = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[45][31].memc__dma__read_data        = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[45][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[45][31].memc__dma__read_ready       = pe_array_inst.pe_inst[45].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 46
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[46][0].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[46][0].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[46][0].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[46][0].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[46][0].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[46][0].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[46][0].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[46][0].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[46][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[46][0].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[46][1].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[46][1].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[46][1].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[46][1].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[46][1].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[46][1].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[46][1].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[46][1].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[46][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[46][1].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[46][2].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[46][2].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[46][2].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[46][2].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[46][2].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[46][2].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[46][2].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[46][2].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[46][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[46][2].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[46][3].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[46][3].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[46][3].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[46][3].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[46][3].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[46][3].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[46][3].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[46][3].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[46][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[46][3].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[46][4].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[46][4].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[46][4].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[46][4].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[46][4].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[46][4].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[46][4].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[46][4].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[46][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[46][4].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[46][5].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[46][5].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[46][5].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[46][5].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[46][5].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[46][5].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[46][5].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[46][5].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[46][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[46][5].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[46][6].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[46][6].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[46][6].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[46][6].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[46][6].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[46][6].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[46][6].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[46][6].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[46][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[46][6].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[46][7].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[46][7].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[46][7].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[46][7].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[46][7].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[46][7].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[46][7].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[46][7].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[46][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[46][7].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[46][8].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[46][8].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[46][8].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[46][8].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[46][8].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[46][8].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[46][8].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[46][8].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[46][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[46][8].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[46][9].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[46][9].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[46][9].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[46][9].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[46][9].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[46][9].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[46][9].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[46][9].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[46][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[46][9].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[46][10].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[46][10].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[46][10].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[46][10].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[46][10].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[46][10].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[46][10].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[46][10].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[46][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[46][10].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[46][11].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[46][11].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[46][11].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[46][11].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[46][11].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[46][11].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[46][11].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[46][11].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[46][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[46][11].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[46][12].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[46][12].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[46][12].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[46][12].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[46][12].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[46][12].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[46][12].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[46][12].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[46][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[46][12].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[46][13].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[46][13].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[46][13].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[46][13].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[46][13].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[46][13].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[46][13].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[46][13].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[46][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[46][13].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[46][14].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[46][14].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[46][14].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[46][14].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[46][14].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[46][14].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[46][14].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[46][14].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[46][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[46][14].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[46][15].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[46][15].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[46][15].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[46][15].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[46][15].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[46][15].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[46][15].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[46][15].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[46][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[46][15].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[46][16].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[46][16].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[46][16].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[46][16].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[46][16].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[46][16].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[46][16].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[46][16].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[46][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[46][16].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[46][17].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[46][17].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[46][17].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[46][17].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[46][17].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[46][17].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[46][17].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[46][17].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[46][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[46][17].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[46][18].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[46][18].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[46][18].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[46][18].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[46][18].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[46][18].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[46][18].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[46][18].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[46][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[46][18].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[46][19].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[46][19].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[46][19].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[46][19].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[46][19].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[46][19].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[46][19].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[46][19].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[46][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[46][19].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[46][20].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[46][20].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[46][20].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[46][20].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[46][20].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[46][20].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[46][20].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[46][20].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[46][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[46][20].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[46][21].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[46][21].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[46][21].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[46][21].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[46][21].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[46][21].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[46][21].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[46][21].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[46][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[46][21].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[46][22].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[46][22].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[46][22].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[46][22].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[46][22].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[46][22].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[46][22].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[46][22].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[46][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[46][22].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[46][23].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[46][23].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[46][23].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[46][23].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[46][23].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[46][23].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[46][23].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[46][23].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[46][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[46][23].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[46][24].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[46][24].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[46][24].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[46][24].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[46][24].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[46][24].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[46][24].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[46][24].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[46][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[46][24].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[46][25].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[46][25].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[46][25].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[46][25].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[46][25].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[46][25].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[46][25].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[46][25].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[46][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[46][25].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[46][26].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[46][26].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[46][26].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[46][26].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[46][26].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[46][26].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[46][26].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[46][26].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[46][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[46][26].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[46][27].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[46][27].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[46][27].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[46][27].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[46][27].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[46][27].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[46][27].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[46][27].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[46][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[46][27].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[46][28].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[46][28].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[46][28].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[46][28].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[46][28].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[46][28].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[46][28].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[46][28].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[46][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[46][28].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[46][29].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[46][29].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[46][29].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[46][29].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[46][29].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[46][29].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[46][29].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[46][29].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[46][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[46][29].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[46][30].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[46][30].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[46][30].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[46][30].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[46][30].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[46][30].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[46][30].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[46][30].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[46][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[46][30].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[46][31].dma__memc__write_valid      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[46][31].dma__memc__write_address    = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[46][31].dma__memc__write_data       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[46][31].dma__memc__read_valid       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[46][31].dma__memc__read_address     = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[46][31].dma__memc__read_pause       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[46][31].memc__dma__write_ready      = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[46][31].memc__dma__read_data        = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[46][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[46][31].memc__dma__read_ready       = pe_array_inst.pe_inst[46].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 47
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[47][0].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[47][0].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[47][0].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[47][0].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[47][0].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[47][0].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[47][0].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[47][0].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[47][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[47][0].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[47][1].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[47][1].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[47][1].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[47][1].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[47][1].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[47][1].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[47][1].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[47][1].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[47][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[47][1].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[47][2].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[47][2].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[47][2].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[47][2].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[47][2].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[47][2].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[47][2].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[47][2].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[47][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[47][2].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[47][3].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[47][3].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[47][3].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[47][3].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[47][3].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[47][3].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[47][3].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[47][3].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[47][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[47][3].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[47][4].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[47][4].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[47][4].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[47][4].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[47][4].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[47][4].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[47][4].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[47][4].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[47][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[47][4].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[47][5].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[47][5].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[47][5].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[47][5].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[47][5].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[47][5].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[47][5].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[47][5].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[47][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[47][5].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[47][6].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[47][6].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[47][6].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[47][6].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[47][6].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[47][6].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[47][6].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[47][6].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[47][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[47][6].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[47][7].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[47][7].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[47][7].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[47][7].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[47][7].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[47][7].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[47][7].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[47][7].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[47][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[47][7].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[47][8].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[47][8].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[47][8].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[47][8].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[47][8].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[47][8].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[47][8].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[47][8].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[47][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[47][8].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[47][9].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[47][9].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[47][9].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[47][9].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[47][9].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[47][9].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[47][9].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[47][9].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[47][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[47][9].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[47][10].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[47][10].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[47][10].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[47][10].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[47][10].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[47][10].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[47][10].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[47][10].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[47][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[47][10].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[47][11].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[47][11].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[47][11].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[47][11].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[47][11].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[47][11].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[47][11].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[47][11].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[47][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[47][11].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[47][12].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[47][12].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[47][12].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[47][12].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[47][12].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[47][12].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[47][12].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[47][12].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[47][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[47][12].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[47][13].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[47][13].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[47][13].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[47][13].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[47][13].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[47][13].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[47][13].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[47][13].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[47][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[47][13].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[47][14].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[47][14].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[47][14].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[47][14].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[47][14].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[47][14].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[47][14].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[47][14].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[47][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[47][14].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[47][15].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[47][15].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[47][15].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[47][15].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[47][15].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[47][15].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[47][15].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[47][15].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[47][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[47][15].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[47][16].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[47][16].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[47][16].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[47][16].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[47][16].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[47][16].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[47][16].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[47][16].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[47][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[47][16].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[47][17].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[47][17].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[47][17].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[47][17].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[47][17].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[47][17].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[47][17].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[47][17].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[47][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[47][17].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[47][18].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[47][18].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[47][18].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[47][18].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[47][18].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[47][18].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[47][18].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[47][18].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[47][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[47][18].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[47][19].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[47][19].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[47][19].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[47][19].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[47][19].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[47][19].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[47][19].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[47][19].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[47][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[47][19].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[47][20].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[47][20].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[47][20].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[47][20].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[47][20].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[47][20].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[47][20].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[47][20].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[47][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[47][20].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[47][21].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[47][21].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[47][21].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[47][21].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[47][21].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[47][21].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[47][21].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[47][21].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[47][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[47][21].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[47][22].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[47][22].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[47][22].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[47][22].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[47][22].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[47][22].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[47][22].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[47][22].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[47][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[47][22].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[47][23].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[47][23].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[47][23].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[47][23].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[47][23].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[47][23].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[47][23].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[47][23].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[47][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[47][23].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[47][24].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[47][24].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[47][24].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[47][24].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[47][24].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[47][24].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[47][24].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[47][24].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[47][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[47][24].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[47][25].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[47][25].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[47][25].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[47][25].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[47][25].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[47][25].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[47][25].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[47][25].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[47][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[47][25].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[47][26].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[47][26].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[47][26].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[47][26].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[47][26].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[47][26].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[47][26].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[47][26].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[47][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[47][26].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[47][27].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[47][27].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[47][27].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[47][27].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[47][27].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[47][27].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[47][27].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[47][27].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[47][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[47][27].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[47][28].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[47][28].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[47][28].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[47][28].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[47][28].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[47][28].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[47][28].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[47][28].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[47][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[47][28].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[47][29].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[47][29].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[47][29].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[47][29].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[47][29].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[47][29].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[47][29].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[47][29].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[47][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[47][29].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[47][30].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[47][30].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[47][30].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[47][30].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[47][30].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[47][30].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[47][30].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[47][30].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[47][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[47][30].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[47][31].dma__memc__write_valid      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[47][31].dma__memc__write_address    = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[47][31].dma__memc__write_data       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[47][31].dma__memc__read_valid       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[47][31].dma__memc__read_address     = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[47][31].dma__memc__read_pause       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[47][31].memc__dma__write_ready      = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[47][31].memc__dma__read_data        = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[47][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[47][31].memc__dma__read_ready       = pe_array_inst.pe_inst[47].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 48
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[48][0].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[48][0].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[48][0].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[48][0].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[48][0].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[48][0].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[48][0].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[48][0].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[48][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[48][0].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[48][1].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[48][1].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[48][1].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[48][1].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[48][1].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[48][1].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[48][1].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[48][1].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[48][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[48][1].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[48][2].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[48][2].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[48][2].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[48][2].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[48][2].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[48][2].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[48][2].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[48][2].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[48][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[48][2].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[48][3].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[48][3].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[48][3].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[48][3].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[48][3].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[48][3].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[48][3].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[48][3].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[48][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[48][3].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[48][4].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[48][4].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[48][4].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[48][4].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[48][4].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[48][4].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[48][4].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[48][4].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[48][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[48][4].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[48][5].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[48][5].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[48][5].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[48][5].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[48][5].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[48][5].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[48][5].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[48][5].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[48][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[48][5].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[48][6].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[48][6].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[48][6].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[48][6].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[48][6].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[48][6].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[48][6].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[48][6].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[48][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[48][6].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[48][7].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[48][7].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[48][7].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[48][7].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[48][7].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[48][7].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[48][7].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[48][7].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[48][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[48][7].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[48][8].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[48][8].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[48][8].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[48][8].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[48][8].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[48][8].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[48][8].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[48][8].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[48][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[48][8].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[48][9].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[48][9].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[48][9].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[48][9].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[48][9].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[48][9].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[48][9].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[48][9].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[48][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[48][9].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[48][10].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[48][10].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[48][10].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[48][10].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[48][10].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[48][10].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[48][10].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[48][10].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[48][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[48][10].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[48][11].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[48][11].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[48][11].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[48][11].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[48][11].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[48][11].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[48][11].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[48][11].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[48][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[48][11].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[48][12].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[48][12].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[48][12].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[48][12].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[48][12].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[48][12].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[48][12].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[48][12].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[48][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[48][12].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[48][13].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[48][13].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[48][13].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[48][13].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[48][13].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[48][13].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[48][13].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[48][13].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[48][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[48][13].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[48][14].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[48][14].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[48][14].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[48][14].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[48][14].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[48][14].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[48][14].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[48][14].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[48][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[48][14].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[48][15].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[48][15].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[48][15].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[48][15].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[48][15].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[48][15].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[48][15].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[48][15].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[48][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[48][15].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[48][16].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[48][16].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[48][16].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[48][16].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[48][16].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[48][16].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[48][16].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[48][16].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[48][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[48][16].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[48][17].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[48][17].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[48][17].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[48][17].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[48][17].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[48][17].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[48][17].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[48][17].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[48][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[48][17].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[48][18].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[48][18].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[48][18].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[48][18].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[48][18].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[48][18].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[48][18].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[48][18].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[48][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[48][18].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[48][19].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[48][19].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[48][19].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[48][19].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[48][19].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[48][19].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[48][19].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[48][19].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[48][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[48][19].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[48][20].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[48][20].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[48][20].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[48][20].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[48][20].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[48][20].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[48][20].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[48][20].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[48][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[48][20].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[48][21].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[48][21].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[48][21].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[48][21].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[48][21].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[48][21].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[48][21].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[48][21].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[48][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[48][21].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[48][22].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[48][22].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[48][22].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[48][22].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[48][22].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[48][22].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[48][22].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[48][22].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[48][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[48][22].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[48][23].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[48][23].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[48][23].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[48][23].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[48][23].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[48][23].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[48][23].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[48][23].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[48][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[48][23].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[48][24].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[48][24].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[48][24].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[48][24].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[48][24].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[48][24].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[48][24].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[48][24].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[48][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[48][24].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[48][25].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[48][25].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[48][25].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[48][25].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[48][25].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[48][25].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[48][25].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[48][25].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[48][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[48][25].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[48][26].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[48][26].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[48][26].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[48][26].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[48][26].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[48][26].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[48][26].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[48][26].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[48][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[48][26].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[48][27].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[48][27].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[48][27].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[48][27].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[48][27].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[48][27].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[48][27].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[48][27].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[48][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[48][27].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[48][28].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[48][28].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[48][28].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[48][28].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[48][28].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[48][28].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[48][28].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[48][28].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[48][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[48][28].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[48][29].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[48][29].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[48][29].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[48][29].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[48][29].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[48][29].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[48][29].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[48][29].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[48][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[48][29].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[48][30].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[48][30].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[48][30].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[48][30].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[48][30].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[48][30].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[48][30].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[48][30].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[48][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[48][30].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[48][31].dma__memc__write_valid      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[48][31].dma__memc__write_address    = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[48][31].dma__memc__write_data       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[48][31].dma__memc__read_valid       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[48][31].dma__memc__read_address     = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[48][31].dma__memc__read_pause       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[48][31].memc__dma__write_ready      = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[48][31].memc__dma__read_data        = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[48][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[48][31].memc__dma__read_ready       = pe_array_inst.pe_inst[48].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 49
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[49][0].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[49][0].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[49][0].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[49][0].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[49][0].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[49][0].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[49][0].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[49][0].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[49][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[49][0].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[49][1].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[49][1].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[49][1].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[49][1].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[49][1].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[49][1].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[49][1].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[49][1].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[49][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[49][1].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[49][2].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[49][2].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[49][2].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[49][2].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[49][2].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[49][2].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[49][2].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[49][2].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[49][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[49][2].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[49][3].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[49][3].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[49][3].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[49][3].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[49][3].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[49][3].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[49][3].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[49][3].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[49][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[49][3].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[49][4].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[49][4].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[49][4].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[49][4].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[49][4].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[49][4].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[49][4].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[49][4].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[49][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[49][4].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[49][5].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[49][5].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[49][5].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[49][5].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[49][5].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[49][5].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[49][5].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[49][5].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[49][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[49][5].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[49][6].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[49][6].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[49][6].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[49][6].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[49][6].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[49][6].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[49][6].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[49][6].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[49][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[49][6].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[49][7].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[49][7].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[49][7].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[49][7].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[49][7].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[49][7].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[49][7].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[49][7].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[49][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[49][7].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[49][8].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[49][8].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[49][8].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[49][8].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[49][8].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[49][8].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[49][8].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[49][8].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[49][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[49][8].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[49][9].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[49][9].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[49][9].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[49][9].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[49][9].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[49][9].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[49][9].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[49][9].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[49][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[49][9].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[49][10].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[49][10].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[49][10].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[49][10].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[49][10].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[49][10].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[49][10].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[49][10].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[49][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[49][10].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[49][11].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[49][11].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[49][11].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[49][11].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[49][11].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[49][11].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[49][11].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[49][11].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[49][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[49][11].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[49][12].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[49][12].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[49][12].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[49][12].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[49][12].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[49][12].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[49][12].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[49][12].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[49][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[49][12].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[49][13].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[49][13].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[49][13].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[49][13].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[49][13].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[49][13].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[49][13].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[49][13].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[49][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[49][13].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[49][14].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[49][14].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[49][14].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[49][14].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[49][14].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[49][14].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[49][14].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[49][14].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[49][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[49][14].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[49][15].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[49][15].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[49][15].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[49][15].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[49][15].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[49][15].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[49][15].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[49][15].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[49][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[49][15].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[49][16].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[49][16].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[49][16].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[49][16].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[49][16].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[49][16].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[49][16].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[49][16].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[49][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[49][16].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[49][17].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[49][17].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[49][17].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[49][17].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[49][17].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[49][17].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[49][17].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[49][17].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[49][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[49][17].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[49][18].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[49][18].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[49][18].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[49][18].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[49][18].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[49][18].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[49][18].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[49][18].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[49][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[49][18].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[49][19].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[49][19].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[49][19].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[49][19].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[49][19].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[49][19].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[49][19].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[49][19].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[49][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[49][19].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[49][20].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[49][20].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[49][20].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[49][20].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[49][20].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[49][20].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[49][20].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[49][20].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[49][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[49][20].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[49][21].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[49][21].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[49][21].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[49][21].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[49][21].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[49][21].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[49][21].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[49][21].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[49][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[49][21].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[49][22].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[49][22].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[49][22].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[49][22].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[49][22].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[49][22].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[49][22].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[49][22].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[49][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[49][22].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[49][23].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[49][23].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[49][23].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[49][23].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[49][23].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[49][23].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[49][23].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[49][23].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[49][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[49][23].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[49][24].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[49][24].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[49][24].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[49][24].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[49][24].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[49][24].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[49][24].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[49][24].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[49][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[49][24].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[49][25].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[49][25].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[49][25].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[49][25].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[49][25].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[49][25].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[49][25].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[49][25].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[49][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[49][25].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[49][26].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[49][26].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[49][26].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[49][26].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[49][26].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[49][26].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[49][26].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[49][26].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[49][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[49][26].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[49][27].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[49][27].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[49][27].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[49][27].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[49][27].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[49][27].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[49][27].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[49][27].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[49][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[49][27].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[49][28].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[49][28].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[49][28].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[49][28].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[49][28].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[49][28].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[49][28].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[49][28].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[49][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[49][28].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[49][29].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[49][29].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[49][29].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[49][29].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[49][29].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[49][29].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[49][29].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[49][29].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[49][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[49][29].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[49][30].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[49][30].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[49][30].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[49][30].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[49][30].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[49][30].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[49][30].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[49][30].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[49][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[49][30].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[49][31].dma__memc__write_valid      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[49][31].dma__memc__write_address    = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[49][31].dma__memc__write_data       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[49][31].dma__memc__read_valid       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[49][31].dma__memc__read_address     = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[49][31].dma__memc__read_pause       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[49][31].memc__dma__write_ready      = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[49][31].memc__dma__read_data        = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[49][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[49][31].memc__dma__read_ready       = pe_array_inst.pe_inst[49].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 50
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[50][0].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[50][0].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[50][0].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[50][0].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[50][0].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[50][0].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[50][0].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[50][0].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[50][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[50][0].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[50][1].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[50][1].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[50][1].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[50][1].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[50][1].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[50][1].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[50][1].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[50][1].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[50][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[50][1].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[50][2].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[50][2].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[50][2].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[50][2].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[50][2].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[50][2].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[50][2].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[50][2].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[50][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[50][2].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[50][3].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[50][3].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[50][3].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[50][3].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[50][3].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[50][3].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[50][3].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[50][3].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[50][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[50][3].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[50][4].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[50][4].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[50][4].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[50][4].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[50][4].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[50][4].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[50][4].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[50][4].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[50][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[50][4].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[50][5].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[50][5].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[50][5].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[50][5].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[50][5].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[50][5].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[50][5].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[50][5].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[50][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[50][5].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[50][6].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[50][6].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[50][6].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[50][6].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[50][6].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[50][6].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[50][6].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[50][6].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[50][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[50][6].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[50][7].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[50][7].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[50][7].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[50][7].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[50][7].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[50][7].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[50][7].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[50][7].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[50][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[50][7].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[50][8].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[50][8].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[50][8].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[50][8].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[50][8].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[50][8].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[50][8].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[50][8].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[50][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[50][8].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[50][9].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[50][9].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[50][9].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[50][9].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[50][9].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[50][9].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[50][9].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[50][9].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[50][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[50][9].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[50][10].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[50][10].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[50][10].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[50][10].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[50][10].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[50][10].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[50][10].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[50][10].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[50][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[50][10].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[50][11].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[50][11].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[50][11].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[50][11].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[50][11].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[50][11].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[50][11].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[50][11].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[50][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[50][11].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[50][12].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[50][12].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[50][12].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[50][12].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[50][12].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[50][12].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[50][12].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[50][12].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[50][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[50][12].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[50][13].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[50][13].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[50][13].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[50][13].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[50][13].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[50][13].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[50][13].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[50][13].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[50][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[50][13].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[50][14].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[50][14].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[50][14].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[50][14].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[50][14].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[50][14].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[50][14].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[50][14].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[50][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[50][14].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[50][15].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[50][15].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[50][15].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[50][15].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[50][15].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[50][15].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[50][15].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[50][15].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[50][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[50][15].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[50][16].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[50][16].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[50][16].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[50][16].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[50][16].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[50][16].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[50][16].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[50][16].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[50][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[50][16].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[50][17].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[50][17].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[50][17].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[50][17].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[50][17].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[50][17].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[50][17].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[50][17].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[50][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[50][17].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[50][18].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[50][18].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[50][18].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[50][18].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[50][18].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[50][18].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[50][18].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[50][18].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[50][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[50][18].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[50][19].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[50][19].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[50][19].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[50][19].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[50][19].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[50][19].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[50][19].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[50][19].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[50][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[50][19].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[50][20].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[50][20].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[50][20].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[50][20].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[50][20].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[50][20].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[50][20].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[50][20].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[50][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[50][20].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[50][21].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[50][21].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[50][21].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[50][21].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[50][21].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[50][21].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[50][21].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[50][21].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[50][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[50][21].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[50][22].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[50][22].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[50][22].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[50][22].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[50][22].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[50][22].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[50][22].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[50][22].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[50][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[50][22].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[50][23].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[50][23].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[50][23].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[50][23].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[50][23].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[50][23].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[50][23].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[50][23].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[50][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[50][23].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[50][24].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[50][24].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[50][24].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[50][24].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[50][24].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[50][24].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[50][24].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[50][24].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[50][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[50][24].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[50][25].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[50][25].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[50][25].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[50][25].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[50][25].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[50][25].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[50][25].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[50][25].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[50][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[50][25].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[50][26].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[50][26].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[50][26].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[50][26].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[50][26].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[50][26].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[50][26].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[50][26].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[50][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[50][26].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[50][27].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[50][27].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[50][27].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[50][27].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[50][27].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[50][27].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[50][27].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[50][27].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[50][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[50][27].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[50][28].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[50][28].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[50][28].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[50][28].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[50][28].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[50][28].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[50][28].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[50][28].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[50][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[50][28].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[50][29].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[50][29].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[50][29].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[50][29].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[50][29].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[50][29].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[50][29].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[50][29].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[50][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[50][29].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[50][30].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[50][30].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[50][30].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[50][30].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[50][30].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[50][30].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[50][30].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[50][30].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[50][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[50][30].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[50][31].dma__memc__write_valid      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[50][31].dma__memc__write_address    = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[50][31].dma__memc__write_data       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[50][31].dma__memc__read_valid       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[50][31].dma__memc__read_address     = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[50][31].dma__memc__read_pause       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[50][31].memc__dma__write_ready      = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[50][31].memc__dma__read_data        = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[50][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[50][31].memc__dma__read_ready       = pe_array_inst.pe_inst[50].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 51
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[51][0].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[51][0].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[51][0].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[51][0].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[51][0].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[51][0].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[51][0].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[51][0].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[51][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[51][0].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[51][1].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[51][1].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[51][1].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[51][1].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[51][1].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[51][1].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[51][1].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[51][1].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[51][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[51][1].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[51][2].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[51][2].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[51][2].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[51][2].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[51][2].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[51][2].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[51][2].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[51][2].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[51][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[51][2].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[51][3].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[51][3].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[51][3].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[51][3].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[51][3].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[51][3].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[51][3].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[51][3].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[51][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[51][3].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[51][4].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[51][4].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[51][4].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[51][4].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[51][4].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[51][4].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[51][4].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[51][4].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[51][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[51][4].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[51][5].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[51][5].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[51][5].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[51][5].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[51][5].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[51][5].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[51][5].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[51][5].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[51][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[51][5].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[51][6].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[51][6].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[51][6].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[51][6].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[51][6].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[51][6].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[51][6].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[51][6].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[51][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[51][6].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[51][7].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[51][7].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[51][7].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[51][7].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[51][7].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[51][7].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[51][7].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[51][7].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[51][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[51][7].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[51][8].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[51][8].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[51][8].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[51][8].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[51][8].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[51][8].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[51][8].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[51][8].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[51][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[51][8].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[51][9].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[51][9].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[51][9].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[51][9].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[51][9].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[51][9].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[51][9].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[51][9].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[51][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[51][9].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[51][10].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[51][10].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[51][10].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[51][10].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[51][10].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[51][10].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[51][10].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[51][10].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[51][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[51][10].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[51][11].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[51][11].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[51][11].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[51][11].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[51][11].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[51][11].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[51][11].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[51][11].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[51][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[51][11].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[51][12].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[51][12].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[51][12].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[51][12].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[51][12].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[51][12].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[51][12].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[51][12].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[51][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[51][12].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[51][13].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[51][13].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[51][13].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[51][13].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[51][13].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[51][13].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[51][13].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[51][13].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[51][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[51][13].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[51][14].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[51][14].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[51][14].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[51][14].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[51][14].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[51][14].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[51][14].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[51][14].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[51][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[51][14].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[51][15].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[51][15].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[51][15].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[51][15].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[51][15].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[51][15].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[51][15].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[51][15].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[51][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[51][15].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[51][16].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[51][16].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[51][16].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[51][16].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[51][16].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[51][16].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[51][16].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[51][16].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[51][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[51][16].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[51][17].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[51][17].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[51][17].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[51][17].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[51][17].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[51][17].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[51][17].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[51][17].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[51][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[51][17].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[51][18].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[51][18].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[51][18].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[51][18].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[51][18].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[51][18].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[51][18].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[51][18].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[51][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[51][18].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[51][19].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[51][19].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[51][19].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[51][19].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[51][19].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[51][19].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[51][19].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[51][19].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[51][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[51][19].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[51][20].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[51][20].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[51][20].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[51][20].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[51][20].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[51][20].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[51][20].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[51][20].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[51][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[51][20].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[51][21].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[51][21].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[51][21].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[51][21].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[51][21].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[51][21].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[51][21].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[51][21].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[51][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[51][21].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[51][22].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[51][22].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[51][22].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[51][22].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[51][22].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[51][22].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[51][22].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[51][22].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[51][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[51][22].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[51][23].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[51][23].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[51][23].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[51][23].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[51][23].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[51][23].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[51][23].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[51][23].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[51][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[51][23].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[51][24].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[51][24].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[51][24].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[51][24].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[51][24].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[51][24].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[51][24].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[51][24].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[51][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[51][24].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[51][25].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[51][25].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[51][25].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[51][25].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[51][25].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[51][25].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[51][25].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[51][25].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[51][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[51][25].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[51][26].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[51][26].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[51][26].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[51][26].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[51][26].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[51][26].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[51][26].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[51][26].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[51][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[51][26].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[51][27].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[51][27].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[51][27].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[51][27].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[51][27].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[51][27].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[51][27].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[51][27].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[51][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[51][27].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[51][28].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[51][28].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[51][28].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[51][28].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[51][28].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[51][28].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[51][28].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[51][28].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[51][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[51][28].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[51][29].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[51][29].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[51][29].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[51][29].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[51][29].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[51][29].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[51][29].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[51][29].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[51][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[51][29].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[51][30].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[51][30].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[51][30].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[51][30].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[51][30].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[51][30].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[51][30].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[51][30].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[51][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[51][30].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[51][31].dma__memc__write_valid      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[51][31].dma__memc__write_address    = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[51][31].dma__memc__write_data       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[51][31].dma__memc__read_valid       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[51][31].dma__memc__read_address     = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[51][31].dma__memc__read_pause       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[51][31].memc__dma__write_ready      = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[51][31].memc__dma__read_data        = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[51][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[51][31].memc__dma__read_ready       = pe_array_inst.pe_inst[51].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 52
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[52][0].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[52][0].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[52][0].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[52][0].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[52][0].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[52][0].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[52][0].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[52][0].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[52][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[52][0].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[52][1].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[52][1].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[52][1].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[52][1].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[52][1].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[52][1].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[52][1].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[52][1].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[52][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[52][1].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[52][2].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[52][2].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[52][2].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[52][2].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[52][2].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[52][2].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[52][2].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[52][2].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[52][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[52][2].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[52][3].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[52][3].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[52][3].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[52][3].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[52][3].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[52][3].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[52][3].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[52][3].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[52][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[52][3].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[52][4].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[52][4].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[52][4].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[52][4].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[52][4].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[52][4].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[52][4].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[52][4].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[52][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[52][4].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[52][5].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[52][5].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[52][5].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[52][5].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[52][5].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[52][5].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[52][5].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[52][5].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[52][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[52][5].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[52][6].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[52][6].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[52][6].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[52][6].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[52][6].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[52][6].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[52][6].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[52][6].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[52][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[52][6].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[52][7].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[52][7].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[52][7].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[52][7].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[52][7].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[52][7].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[52][7].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[52][7].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[52][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[52][7].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[52][8].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[52][8].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[52][8].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[52][8].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[52][8].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[52][8].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[52][8].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[52][8].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[52][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[52][8].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[52][9].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[52][9].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[52][9].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[52][9].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[52][9].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[52][9].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[52][9].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[52][9].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[52][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[52][9].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[52][10].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[52][10].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[52][10].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[52][10].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[52][10].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[52][10].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[52][10].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[52][10].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[52][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[52][10].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[52][11].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[52][11].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[52][11].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[52][11].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[52][11].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[52][11].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[52][11].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[52][11].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[52][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[52][11].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[52][12].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[52][12].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[52][12].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[52][12].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[52][12].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[52][12].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[52][12].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[52][12].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[52][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[52][12].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[52][13].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[52][13].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[52][13].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[52][13].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[52][13].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[52][13].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[52][13].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[52][13].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[52][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[52][13].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[52][14].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[52][14].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[52][14].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[52][14].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[52][14].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[52][14].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[52][14].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[52][14].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[52][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[52][14].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[52][15].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[52][15].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[52][15].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[52][15].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[52][15].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[52][15].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[52][15].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[52][15].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[52][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[52][15].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[52][16].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[52][16].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[52][16].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[52][16].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[52][16].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[52][16].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[52][16].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[52][16].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[52][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[52][16].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[52][17].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[52][17].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[52][17].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[52][17].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[52][17].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[52][17].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[52][17].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[52][17].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[52][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[52][17].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[52][18].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[52][18].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[52][18].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[52][18].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[52][18].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[52][18].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[52][18].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[52][18].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[52][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[52][18].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[52][19].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[52][19].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[52][19].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[52][19].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[52][19].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[52][19].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[52][19].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[52][19].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[52][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[52][19].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[52][20].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[52][20].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[52][20].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[52][20].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[52][20].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[52][20].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[52][20].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[52][20].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[52][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[52][20].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[52][21].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[52][21].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[52][21].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[52][21].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[52][21].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[52][21].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[52][21].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[52][21].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[52][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[52][21].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[52][22].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[52][22].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[52][22].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[52][22].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[52][22].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[52][22].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[52][22].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[52][22].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[52][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[52][22].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[52][23].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[52][23].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[52][23].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[52][23].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[52][23].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[52][23].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[52][23].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[52][23].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[52][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[52][23].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[52][24].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[52][24].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[52][24].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[52][24].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[52][24].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[52][24].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[52][24].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[52][24].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[52][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[52][24].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[52][25].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[52][25].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[52][25].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[52][25].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[52][25].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[52][25].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[52][25].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[52][25].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[52][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[52][25].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[52][26].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[52][26].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[52][26].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[52][26].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[52][26].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[52][26].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[52][26].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[52][26].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[52][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[52][26].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[52][27].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[52][27].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[52][27].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[52][27].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[52][27].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[52][27].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[52][27].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[52][27].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[52][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[52][27].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[52][28].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[52][28].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[52][28].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[52][28].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[52][28].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[52][28].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[52][28].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[52][28].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[52][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[52][28].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[52][29].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[52][29].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[52][29].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[52][29].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[52][29].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[52][29].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[52][29].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[52][29].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[52][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[52][29].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[52][30].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[52][30].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[52][30].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[52][30].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[52][30].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[52][30].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[52][30].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[52][30].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[52][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[52][30].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[52][31].dma__memc__write_valid      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[52][31].dma__memc__write_address    = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[52][31].dma__memc__write_data       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[52][31].dma__memc__read_valid       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[52][31].dma__memc__read_address     = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[52][31].dma__memc__read_pause       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[52][31].memc__dma__write_ready      = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[52][31].memc__dma__read_data        = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[52][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[52][31].memc__dma__read_ready       = pe_array_inst.pe_inst[52].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 53
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[53][0].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[53][0].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[53][0].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[53][0].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[53][0].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[53][0].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[53][0].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[53][0].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[53][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[53][0].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[53][1].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[53][1].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[53][1].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[53][1].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[53][1].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[53][1].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[53][1].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[53][1].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[53][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[53][1].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[53][2].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[53][2].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[53][2].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[53][2].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[53][2].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[53][2].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[53][2].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[53][2].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[53][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[53][2].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[53][3].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[53][3].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[53][3].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[53][3].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[53][3].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[53][3].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[53][3].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[53][3].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[53][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[53][3].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[53][4].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[53][4].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[53][4].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[53][4].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[53][4].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[53][4].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[53][4].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[53][4].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[53][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[53][4].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[53][5].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[53][5].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[53][5].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[53][5].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[53][5].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[53][5].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[53][5].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[53][5].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[53][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[53][5].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[53][6].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[53][6].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[53][6].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[53][6].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[53][6].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[53][6].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[53][6].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[53][6].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[53][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[53][6].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[53][7].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[53][7].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[53][7].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[53][7].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[53][7].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[53][7].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[53][7].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[53][7].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[53][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[53][7].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[53][8].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[53][8].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[53][8].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[53][8].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[53][8].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[53][8].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[53][8].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[53][8].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[53][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[53][8].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[53][9].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[53][9].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[53][9].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[53][9].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[53][9].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[53][9].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[53][9].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[53][9].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[53][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[53][9].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[53][10].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[53][10].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[53][10].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[53][10].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[53][10].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[53][10].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[53][10].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[53][10].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[53][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[53][10].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[53][11].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[53][11].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[53][11].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[53][11].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[53][11].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[53][11].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[53][11].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[53][11].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[53][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[53][11].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[53][12].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[53][12].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[53][12].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[53][12].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[53][12].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[53][12].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[53][12].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[53][12].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[53][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[53][12].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[53][13].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[53][13].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[53][13].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[53][13].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[53][13].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[53][13].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[53][13].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[53][13].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[53][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[53][13].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[53][14].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[53][14].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[53][14].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[53][14].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[53][14].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[53][14].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[53][14].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[53][14].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[53][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[53][14].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[53][15].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[53][15].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[53][15].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[53][15].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[53][15].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[53][15].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[53][15].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[53][15].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[53][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[53][15].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[53][16].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[53][16].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[53][16].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[53][16].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[53][16].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[53][16].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[53][16].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[53][16].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[53][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[53][16].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[53][17].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[53][17].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[53][17].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[53][17].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[53][17].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[53][17].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[53][17].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[53][17].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[53][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[53][17].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[53][18].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[53][18].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[53][18].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[53][18].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[53][18].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[53][18].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[53][18].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[53][18].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[53][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[53][18].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[53][19].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[53][19].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[53][19].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[53][19].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[53][19].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[53][19].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[53][19].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[53][19].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[53][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[53][19].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[53][20].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[53][20].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[53][20].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[53][20].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[53][20].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[53][20].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[53][20].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[53][20].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[53][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[53][20].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[53][21].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[53][21].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[53][21].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[53][21].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[53][21].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[53][21].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[53][21].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[53][21].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[53][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[53][21].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[53][22].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[53][22].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[53][22].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[53][22].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[53][22].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[53][22].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[53][22].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[53][22].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[53][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[53][22].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[53][23].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[53][23].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[53][23].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[53][23].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[53][23].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[53][23].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[53][23].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[53][23].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[53][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[53][23].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[53][24].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[53][24].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[53][24].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[53][24].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[53][24].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[53][24].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[53][24].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[53][24].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[53][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[53][24].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[53][25].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[53][25].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[53][25].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[53][25].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[53][25].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[53][25].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[53][25].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[53][25].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[53][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[53][25].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[53][26].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[53][26].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[53][26].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[53][26].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[53][26].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[53][26].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[53][26].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[53][26].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[53][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[53][26].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[53][27].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[53][27].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[53][27].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[53][27].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[53][27].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[53][27].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[53][27].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[53][27].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[53][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[53][27].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[53][28].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[53][28].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[53][28].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[53][28].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[53][28].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[53][28].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[53][28].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[53][28].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[53][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[53][28].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[53][29].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[53][29].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[53][29].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[53][29].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[53][29].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[53][29].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[53][29].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[53][29].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[53][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[53][29].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[53][30].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[53][30].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[53][30].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[53][30].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[53][30].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[53][30].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[53][30].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[53][30].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[53][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[53][30].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[53][31].dma__memc__write_valid      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[53][31].dma__memc__write_address    = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[53][31].dma__memc__write_data       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[53][31].dma__memc__read_valid       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[53][31].dma__memc__read_address     = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[53][31].dma__memc__read_pause       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[53][31].memc__dma__write_ready      = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[53][31].memc__dma__read_data        = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[53][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[53][31].memc__dma__read_ready       = pe_array_inst.pe_inst[53].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 54
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[54][0].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[54][0].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[54][0].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[54][0].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[54][0].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[54][0].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[54][0].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[54][0].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[54][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[54][0].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[54][1].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[54][1].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[54][1].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[54][1].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[54][1].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[54][1].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[54][1].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[54][1].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[54][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[54][1].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[54][2].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[54][2].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[54][2].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[54][2].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[54][2].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[54][2].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[54][2].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[54][2].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[54][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[54][2].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[54][3].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[54][3].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[54][3].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[54][3].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[54][3].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[54][3].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[54][3].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[54][3].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[54][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[54][3].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[54][4].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[54][4].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[54][4].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[54][4].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[54][4].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[54][4].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[54][4].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[54][4].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[54][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[54][4].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[54][5].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[54][5].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[54][5].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[54][5].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[54][5].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[54][5].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[54][5].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[54][5].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[54][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[54][5].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[54][6].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[54][6].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[54][6].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[54][6].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[54][6].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[54][6].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[54][6].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[54][6].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[54][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[54][6].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[54][7].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[54][7].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[54][7].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[54][7].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[54][7].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[54][7].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[54][7].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[54][7].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[54][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[54][7].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[54][8].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[54][8].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[54][8].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[54][8].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[54][8].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[54][8].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[54][8].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[54][8].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[54][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[54][8].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[54][9].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[54][9].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[54][9].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[54][9].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[54][9].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[54][9].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[54][9].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[54][9].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[54][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[54][9].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[54][10].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[54][10].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[54][10].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[54][10].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[54][10].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[54][10].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[54][10].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[54][10].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[54][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[54][10].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[54][11].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[54][11].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[54][11].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[54][11].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[54][11].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[54][11].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[54][11].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[54][11].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[54][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[54][11].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[54][12].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[54][12].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[54][12].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[54][12].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[54][12].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[54][12].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[54][12].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[54][12].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[54][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[54][12].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[54][13].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[54][13].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[54][13].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[54][13].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[54][13].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[54][13].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[54][13].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[54][13].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[54][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[54][13].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[54][14].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[54][14].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[54][14].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[54][14].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[54][14].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[54][14].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[54][14].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[54][14].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[54][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[54][14].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[54][15].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[54][15].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[54][15].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[54][15].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[54][15].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[54][15].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[54][15].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[54][15].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[54][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[54][15].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[54][16].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[54][16].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[54][16].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[54][16].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[54][16].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[54][16].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[54][16].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[54][16].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[54][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[54][16].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[54][17].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[54][17].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[54][17].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[54][17].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[54][17].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[54][17].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[54][17].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[54][17].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[54][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[54][17].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[54][18].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[54][18].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[54][18].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[54][18].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[54][18].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[54][18].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[54][18].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[54][18].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[54][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[54][18].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[54][19].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[54][19].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[54][19].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[54][19].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[54][19].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[54][19].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[54][19].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[54][19].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[54][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[54][19].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[54][20].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[54][20].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[54][20].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[54][20].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[54][20].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[54][20].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[54][20].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[54][20].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[54][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[54][20].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[54][21].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[54][21].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[54][21].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[54][21].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[54][21].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[54][21].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[54][21].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[54][21].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[54][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[54][21].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[54][22].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[54][22].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[54][22].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[54][22].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[54][22].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[54][22].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[54][22].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[54][22].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[54][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[54][22].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[54][23].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[54][23].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[54][23].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[54][23].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[54][23].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[54][23].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[54][23].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[54][23].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[54][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[54][23].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[54][24].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[54][24].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[54][24].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[54][24].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[54][24].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[54][24].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[54][24].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[54][24].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[54][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[54][24].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[54][25].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[54][25].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[54][25].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[54][25].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[54][25].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[54][25].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[54][25].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[54][25].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[54][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[54][25].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[54][26].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[54][26].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[54][26].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[54][26].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[54][26].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[54][26].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[54][26].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[54][26].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[54][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[54][26].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[54][27].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[54][27].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[54][27].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[54][27].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[54][27].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[54][27].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[54][27].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[54][27].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[54][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[54][27].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[54][28].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[54][28].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[54][28].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[54][28].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[54][28].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[54][28].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[54][28].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[54][28].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[54][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[54][28].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[54][29].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[54][29].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[54][29].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[54][29].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[54][29].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[54][29].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[54][29].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[54][29].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[54][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[54][29].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[54][30].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[54][30].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[54][30].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[54][30].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[54][30].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[54][30].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[54][30].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[54][30].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[54][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[54][30].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[54][31].dma__memc__write_valid      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[54][31].dma__memc__write_address    = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[54][31].dma__memc__write_data       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[54][31].dma__memc__read_valid       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[54][31].dma__memc__read_address     = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[54][31].dma__memc__read_pause       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[54][31].memc__dma__write_ready      = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[54][31].memc__dma__read_data        = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[54][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[54][31].memc__dma__read_ready       = pe_array_inst.pe_inst[54].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 55
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[55][0].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[55][0].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[55][0].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[55][0].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[55][0].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[55][0].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[55][0].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[55][0].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[55][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[55][0].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[55][1].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[55][1].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[55][1].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[55][1].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[55][1].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[55][1].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[55][1].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[55][1].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[55][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[55][1].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[55][2].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[55][2].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[55][2].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[55][2].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[55][2].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[55][2].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[55][2].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[55][2].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[55][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[55][2].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[55][3].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[55][3].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[55][3].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[55][3].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[55][3].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[55][3].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[55][3].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[55][3].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[55][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[55][3].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[55][4].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[55][4].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[55][4].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[55][4].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[55][4].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[55][4].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[55][4].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[55][4].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[55][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[55][4].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[55][5].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[55][5].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[55][5].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[55][5].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[55][5].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[55][5].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[55][5].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[55][5].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[55][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[55][5].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[55][6].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[55][6].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[55][6].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[55][6].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[55][6].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[55][6].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[55][6].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[55][6].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[55][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[55][6].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[55][7].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[55][7].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[55][7].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[55][7].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[55][7].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[55][7].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[55][7].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[55][7].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[55][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[55][7].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[55][8].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[55][8].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[55][8].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[55][8].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[55][8].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[55][8].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[55][8].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[55][8].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[55][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[55][8].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[55][9].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[55][9].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[55][9].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[55][9].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[55][9].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[55][9].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[55][9].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[55][9].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[55][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[55][9].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[55][10].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[55][10].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[55][10].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[55][10].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[55][10].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[55][10].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[55][10].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[55][10].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[55][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[55][10].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[55][11].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[55][11].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[55][11].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[55][11].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[55][11].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[55][11].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[55][11].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[55][11].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[55][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[55][11].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[55][12].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[55][12].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[55][12].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[55][12].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[55][12].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[55][12].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[55][12].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[55][12].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[55][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[55][12].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[55][13].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[55][13].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[55][13].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[55][13].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[55][13].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[55][13].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[55][13].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[55][13].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[55][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[55][13].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[55][14].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[55][14].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[55][14].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[55][14].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[55][14].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[55][14].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[55][14].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[55][14].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[55][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[55][14].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[55][15].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[55][15].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[55][15].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[55][15].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[55][15].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[55][15].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[55][15].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[55][15].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[55][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[55][15].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[55][16].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[55][16].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[55][16].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[55][16].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[55][16].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[55][16].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[55][16].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[55][16].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[55][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[55][16].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[55][17].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[55][17].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[55][17].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[55][17].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[55][17].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[55][17].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[55][17].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[55][17].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[55][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[55][17].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[55][18].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[55][18].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[55][18].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[55][18].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[55][18].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[55][18].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[55][18].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[55][18].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[55][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[55][18].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[55][19].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[55][19].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[55][19].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[55][19].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[55][19].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[55][19].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[55][19].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[55][19].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[55][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[55][19].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[55][20].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[55][20].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[55][20].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[55][20].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[55][20].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[55][20].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[55][20].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[55][20].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[55][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[55][20].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[55][21].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[55][21].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[55][21].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[55][21].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[55][21].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[55][21].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[55][21].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[55][21].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[55][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[55][21].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[55][22].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[55][22].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[55][22].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[55][22].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[55][22].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[55][22].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[55][22].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[55][22].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[55][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[55][22].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[55][23].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[55][23].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[55][23].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[55][23].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[55][23].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[55][23].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[55][23].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[55][23].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[55][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[55][23].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[55][24].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[55][24].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[55][24].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[55][24].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[55][24].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[55][24].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[55][24].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[55][24].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[55][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[55][24].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[55][25].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[55][25].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[55][25].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[55][25].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[55][25].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[55][25].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[55][25].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[55][25].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[55][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[55][25].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[55][26].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[55][26].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[55][26].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[55][26].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[55][26].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[55][26].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[55][26].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[55][26].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[55][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[55][26].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[55][27].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[55][27].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[55][27].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[55][27].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[55][27].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[55][27].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[55][27].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[55][27].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[55][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[55][27].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[55][28].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[55][28].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[55][28].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[55][28].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[55][28].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[55][28].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[55][28].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[55][28].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[55][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[55][28].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[55][29].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[55][29].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[55][29].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[55][29].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[55][29].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[55][29].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[55][29].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[55][29].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[55][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[55][29].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[55][30].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[55][30].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[55][30].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[55][30].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[55][30].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[55][30].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[55][30].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[55][30].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[55][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[55][30].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[55][31].dma__memc__write_valid      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[55][31].dma__memc__write_address    = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[55][31].dma__memc__write_data       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[55][31].dma__memc__read_valid       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[55][31].dma__memc__read_address     = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[55][31].dma__memc__read_pause       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[55][31].memc__dma__write_ready      = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[55][31].memc__dma__read_data        = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[55][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[55][31].memc__dma__read_ready       = pe_array_inst.pe_inst[55].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 56
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[56][0].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[56][0].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[56][0].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[56][0].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[56][0].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[56][0].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[56][0].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[56][0].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[56][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[56][0].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[56][1].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[56][1].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[56][1].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[56][1].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[56][1].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[56][1].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[56][1].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[56][1].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[56][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[56][1].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[56][2].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[56][2].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[56][2].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[56][2].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[56][2].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[56][2].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[56][2].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[56][2].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[56][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[56][2].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[56][3].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[56][3].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[56][3].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[56][3].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[56][3].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[56][3].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[56][3].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[56][3].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[56][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[56][3].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[56][4].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[56][4].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[56][4].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[56][4].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[56][4].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[56][4].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[56][4].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[56][4].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[56][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[56][4].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[56][5].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[56][5].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[56][5].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[56][5].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[56][5].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[56][5].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[56][5].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[56][5].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[56][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[56][5].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[56][6].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[56][6].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[56][6].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[56][6].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[56][6].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[56][6].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[56][6].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[56][6].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[56][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[56][6].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[56][7].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[56][7].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[56][7].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[56][7].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[56][7].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[56][7].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[56][7].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[56][7].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[56][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[56][7].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[56][8].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[56][8].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[56][8].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[56][8].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[56][8].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[56][8].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[56][8].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[56][8].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[56][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[56][8].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[56][9].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[56][9].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[56][9].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[56][9].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[56][9].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[56][9].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[56][9].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[56][9].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[56][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[56][9].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[56][10].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[56][10].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[56][10].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[56][10].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[56][10].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[56][10].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[56][10].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[56][10].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[56][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[56][10].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[56][11].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[56][11].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[56][11].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[56][11].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[56][11].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[56][11].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[56][11].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[56][11].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[56][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[56][11].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[56][12].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[56][12].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[56][12].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[56][12].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[56][12].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[56][12].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[56][12].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[56][12].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[56][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[56][12].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[56][13].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[56][13].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[56][13].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[56][13].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[56][13].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[56][13].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[56][13].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[56][13].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[56][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[56][13].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[56][14].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[56][14].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[56][14].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[56][14].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[56][14].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[56][14].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[56][14].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[56][14].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[56][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[56][14].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[56][15].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[56][15].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[56][15].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[56][15].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[56][15].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[56][15].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[56][15].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[56][15].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[56][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[56][15].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[56][16].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[56][16].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[56][16].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[56][16].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[56][16].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[56][16].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[56][16].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[56][16].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[56][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[56][16].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[56][17].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[56][17].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[56][17].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[56][17].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[56][17].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[56][17].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[56][17].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[56][17].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[56][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[56][17].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[56][18].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[56][18].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[56][18].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[56][18].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[56][18].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[56][18].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[56][18].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[56][18].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[56][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[56][18].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[56][19].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[56][19].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[56][19].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[56][19].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[56][19].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[56][19].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[56][19].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[56][19].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[56][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[56][19].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[56][20].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[56][20].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[56][20].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[56][20].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[56][20].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[56][20].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[56][20].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[56][20].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[56][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[56][20].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[56][21].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[56][21].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[56][21].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[56][21].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[56][21].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[56][21].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[56][21].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[56][21].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[56][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[56][21].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[56][22].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[56][22].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[56][22].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[56][22].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[56][22].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[56][22].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[56][22].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[56][22].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[56][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[56][22].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[56][23].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[56][23].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[56][23].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[56][23].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[56][23].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[56][23].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[56][23].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[56][23].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[56][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[56][23].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[56][24].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[56][24].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[56][24].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[56][24].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[56][24].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[56][24].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[56][24].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[56][24].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[56][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[56][24].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[56][25].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[56][25].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[56][25].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[56][25].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[56][25].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[56][25].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[56][25].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[56][25].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[56][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[56][25].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[56][26].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[56][26].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[56][26].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[56][26].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[56][26].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[56][26].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[56][26].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[56][26].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[56][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[56][26].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[56][27].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[56][27].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[56][27].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[56][27].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[56][27].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[56][27].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[56][27].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[56][27].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[56][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[56][27].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[56][28].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[56][28].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[56][28].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[56][28].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[56][28].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[56][28].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[56][28].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[56][28].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[56][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[56][28].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[56][29].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[56][29].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[56][29].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[56][29].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[56][29].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[56][29].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[56][29].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[56][29].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[56][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[56][29].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[56][30].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[56][30].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[56][30].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[56][30].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[56][30].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[56][30].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[56][30].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[56][30].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[56][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[56][30].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[56][31].dma__memc__write_valid      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[56][31].dma__memc__write_address    = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[56][31].dma__memc__write_data       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[56][31].dma__memc__read_valid       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[56][31].dma__memc__read_address     = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[56][31].dma__memc__read_pause       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[56][31].memc__dma__write_ready      = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[56][31].memc__dma__read_data        = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[56][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[56][31].memc__dma__read_ready       = pe_array_inst.pe_inst[56].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 57
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[57][0].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[57][0].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[57][0].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[57][0].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[57][0].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[57][0].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[57][0].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[57][0].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[57][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[57][0].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[57][1].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[57][1].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[57][1].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[57][1].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[57][1].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[57][1].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[57][1].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[57][1].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[57][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[57][1].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[57][2].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[57][2].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[57][2].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[57][2].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[57][2].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[57][2].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[57][2].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[57][2].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[57][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[57][2].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[57][3].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[57][3].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[57][3].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[57][3].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[57][3].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[57][3].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[57][3].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[57][3].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[57][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[57][3].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[57][4].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[57][4].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[57][4].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[57][4].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[57][4].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[57][4].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[57][4].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[57][4].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[57][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[57][4].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[57][5].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[57][5].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[57][5].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[57][5].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[57][5].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[57][5].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[57][5].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[57][5].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[57][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[57][5].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[57][6].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[57][6].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[57][6].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[57][6].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[57][6].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[57][6].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[57][6].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[57][6].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[57][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[57][6].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[57][7].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[57][7].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[57][7].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[57][7].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[57][7].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[57][7].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[57][7].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[57][7].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[57][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[57][7].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[57][8].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[57][8].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[57][8].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[57][8].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[57][8].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[57][8].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[57][8].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[57][8].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[57][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[57][8].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[57][9].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[57][9].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[57][9].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[57][9].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[57][9].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[57][9].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[57][9].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[57][9].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[57][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[57][9].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[57][10].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[57][10].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[57][10].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[57][10].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[57][10].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[57][10].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[57][10].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[57][10].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[57][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[57][10].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[57][11].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[57][11].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[57][11].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[57][11].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[57][11].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[57][11].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[57][11].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[57][11].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[57][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[57][11].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[57][12].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[57][12].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[57][12].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[57][12].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[57][12].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[57][12].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[57][12].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[57][12].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[57][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[57][12].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[57][13].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[57][13].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[57][13].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[57][13].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[57][13].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[57][13].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[57][13].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[57][13].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[57][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[57][13].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[57][14].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[57][14].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[57][14].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[57][14].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[57][14].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[57][14].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[57][14].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[57][14].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[57][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[57][14].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[57][15].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[57][15].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[57][15].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[57][15].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[57][15].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[57][15].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[57][15].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[57][15].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[57][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[57][15].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[57][16].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[57][16].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[57][16].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[57][16].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[57][16].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[57][16].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[57][16].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[57][16].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[57][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[57][16].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[57][17].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[57][17].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[57][17].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[57][17].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[57][17].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[57][17].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[57][17].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[57][17].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[57][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[57][17].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[57][18].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[57][18].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[57][18].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[57][18].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[57][18].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[57][18].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[57][18].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[57][18].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[57][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[57][18].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[57][19].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[57][19].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[57][19].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[57][19].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[57][19].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[57][19].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[57][19].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[57][19].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[57][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[57][19].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[57][20].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[57][20].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[57][20].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[57][20].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[57][20].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[57][20].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[57][20].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[57][20].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[57][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[57][20].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[57][21].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[57][21].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[57][21].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[57][21].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[57][21].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[57][21].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[57][21].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[57][21].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[57][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[57][21].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[57][22].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[57][22].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[57][22].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[57][22].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[57][22].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[57][22].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[57][22].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[57][22].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[57][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[57][22].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[57][23].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[57][23].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[57][23].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[57][23].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[57][23].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[57][23].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[57][23].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[57][23].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[57][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[57][23].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[57][24].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[57][24].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[57][24].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[57][24].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[57][24].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[57][24].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[57][24].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[57][24].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[57][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[57][24].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[57][25].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[57][25].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[57][25].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[57][25].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[57][25].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[57][25].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[57][25].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[57][25].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[57][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[57][25].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[57][26].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[57][26].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[57][26].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[57][26].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[57][26].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[57][26].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[57][26].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[57][26].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[57][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[57][26].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[57][27].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[57][27].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[57][27].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[57][27].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[57][27].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[57][27].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[57][27].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[57][27].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[57][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[57][27].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[57][28].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[57][28].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[57][28].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[57][28].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[57][28].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[57][28].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[57][28].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[57][28].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[57][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[57][28].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[57][29].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[57][29].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[57][29].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[57][29].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[57][29].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[57][29].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[57][29].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[57][29].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[57][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[57][29].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[57][30].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[57][30].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[57][30].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[57][30].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[57][30].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[57][30].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[57][30].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[57][30].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[57][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[57][30].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[57][31].dma__memc__write_valid      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[57][31].dma__memc__write_address    = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[57][31].dma__memc__write_data       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[57][31].dma__memc__read_valid       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[57][31].dma__memc__read_address     = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[57][31].dma__memc__read_pause       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[57][31].memc__dma__write_ready      = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[57][31].memc__dma__read_data        = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[57][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[57][31].memc__dma__read_ready       = pe_array_inst.pe_inst[57].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 58
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[58][0].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[58][0].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[58][0].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[58][0].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[58][0].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[58][0].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[58][0].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[58][0].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[58][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[58][0].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[58][1].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[58][1].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[58][1].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[58][1].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[58][1].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[58][1].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[58][1].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[58][1].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[58][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[58][1].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[58][2].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[58][2].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[58][2].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[58][2].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[58][2].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[58][2].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[58][2].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[58][2].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[58][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[58][2].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[58][3].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[58][3].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[58][3].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[58][3].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[58][3].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[58][3].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[58][3].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[58][3].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[58][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[58][3].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[58][4].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[58][4].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[58][4].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[58][4].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[58][4].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[58][4].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[58][4].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[58][4].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[58][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[58][4].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[58][5].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[58][5].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[58][5].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[58][5].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[58][5].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[58][5].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[58][5].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[58][5].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[58][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[58][5].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[58][6].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[58][6].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[58][6].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[58][6].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[58][6].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[58][6].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[58][6].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[58][6].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[58][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[58][6].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[58][7].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[58][7].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[58][7].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[58][7].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[58][7].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[58][7].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[58][7].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[58][7].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[58][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[58][7].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[58][8].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[58][8].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[58][8].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[58][8].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[58][8].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[58][8].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[58][8].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[58][8].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[58][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[58][8].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[58][9].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[58][9].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[58][9].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[58][9].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[58][9].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[58][9].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[58][9].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[58][9].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[58][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[58][9].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[58][10].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[58][10].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[58][10].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[58][10].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[58][10].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[58][10].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[58][10].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[58][10].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[58][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[58][10].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[58][11].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[58][11].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[58][11].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[58][11].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[58][11].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[58][11].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[58][11].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[58][11].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[58][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[58][11].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[58][12].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[58][12].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[58][12].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[58][12].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[58][12].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[58][12].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[58][12].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[58][12].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[58][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[58][12].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[58][13].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[58][13].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[58][13].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[58][13].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[58][13].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[58][13].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[58][13].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[58][13].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[58][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[58][13].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[58][14].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[58][14].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[58][14].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[58][14].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[58][14].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[58][14].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[58][14].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[58][14].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[58][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[58][14].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[58][15].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[58][15].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[58][15].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[58][15].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[58][15].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[58][15].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[58][15].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[58][15].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[58][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[58][15].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[58][16].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[58][16].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[58][16].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[58][16].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[58][16].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[58][16].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[58][16].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[58][16].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[58][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[58][16].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[58][17].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[58][17].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[58][17].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[58][17].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[58][17].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[58][17].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[58][17].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[58][17].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[58][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[58][17].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[58][18].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[58][18].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[58][18].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[58][18].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[58][18].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[58][18].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[58][18].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[58][18].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[58][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[58][18].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[58][19].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[58][19].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[58][19].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[58][19].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[58][19].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[58][19].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[58][19].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[58][19].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[58][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[58][19].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[58][20].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[58][20].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[58][20].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[58][20].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[58][20].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[58][20].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[58][20].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[58][20].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[58][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[58][20].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[58][21].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[58][21].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[58][21].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[58][21].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[58][21].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[58][21].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[58][21].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[58][21].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[58][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[58][21].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[58][22].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[58][22].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[58][22].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[58][22].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[58][22].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[58][22].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[58][22].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[58][22].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[58][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[58][22].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[58][23].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[58][23].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[58][23].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[58][23].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[58][23].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[58][23].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[58][23].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[58][23].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[58][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[58][23].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[58][24].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[58][24].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[58][24].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[58][24].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[58][24].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[58][24].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[58][24].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[58][24].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[58][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[58][24].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[58][25].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[58][25].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[58][25].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[58][25].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[58][25].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[58][25].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[58][25].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[58][25].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[58][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[58][25].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[58][26].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[58][26].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[58][26].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[58][26].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[58][26].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[58][26].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[58][26].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[58][26].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[58][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[58][26].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[58][27].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[58][27].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[58][27].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[58][27].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[58][27].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[58][27].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[58][27].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[58][27].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[58][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[58][27].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[58][28].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[58][28].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[58][28].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[58][28].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[58][28].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[58][28].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[58][28].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[58][28].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[58][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[58][28].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[58][29].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[58][29].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[58][29].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[58][29].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[58][29].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[58][29].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[58][29].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[58][29].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[58][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[58][29].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[58][30].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[58][30].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[58][30].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[58][30].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[58][30].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[58][30].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[58][30].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[58][30].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[58][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[58][30].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[58][31].dma__memc__write_valid      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[58][31].dma__memc__write_address    = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[58][31].dma__memc__write_data       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[58][31].dma__memc__read_valid       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[58][31].dma__memc__read_address     = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[58][31].dma__memc__read_pause       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[58][31].memc__dma__write_ready      = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[58][31].memc__dma__read_data        = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[58][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[58][31].memc__dma__read_ready       = pe_array_inst.pe_inst[58].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 59
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[59][0].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[59][0].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[59][0].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[59][0].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[59][0].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[59][0].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[59][0].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[59][0].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[59][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[59][0].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[59][1].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[59][1].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[59][1].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[59][1].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[59][1].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[59][1].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[59][1].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[59][1].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[59][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[59][1].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[59][2].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[59][2].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[59][2].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[59][2].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[59][2].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[59][2].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[59][2].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[59][2].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[59][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[59][2].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[59][3].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[59][3].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[59][3].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[59][3].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[59][3].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[59][3].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[59][3].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[59][3].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[59][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[59][3].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[59][4].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[59][4].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[59][4].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[59][4].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[59][4].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[59][4].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[59][4].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[59][4].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[59][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[59][4].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[59][5].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[59][5].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[59][5].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[59][5].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[59][5].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[59][5].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[59][5].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[59][5].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[59][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[59][5].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[59][6].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[59][6].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[59][6].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[59][6].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[59][6].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[59][6].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[59][6].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[59][6].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[59][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[59][6].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[59][7].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[59][7].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[59][7].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[59][7].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[59][7].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[59][7].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[59][7].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[59][7].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[59][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[59][7].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[59][8].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[59][8].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[59][8].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[59][8].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[59][8].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[59][8].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[59][8].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[59][8].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[59][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[59][8].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[59][9].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[59][9].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[59][9].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[59][9].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[59][9].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[59][9].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[59][9].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[59][9].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[59][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[59][9].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[59][10].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[59][10].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[59][10].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[59][10].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[59][10].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[59][10].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[59][10].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[59][10].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[59][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[59][10].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[59][11].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[59][11].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[59][11].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[59][11].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[59][11].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[59][11].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[59][11].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[59][11].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[59][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[59][11].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[59][12].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[59][12].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[59][12].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[59][12].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[59][12].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[59][12].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[59][12].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[59][12].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[59][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[59][12].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[59][13].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[59][13].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[59][13].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[59][13].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[59][13].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[59][13].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[59][13].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[59][13].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[59][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[59][13].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[59][14].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[59][14].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[59][14].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[59][14].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[59][14].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[59][14].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[59][14].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[59][14].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[59][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[59][14].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[59][15].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[59][15].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[59][15].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[59][15].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[59][15].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[59][15].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[59][15].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[59][15].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[59][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[59][15].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[59][16].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[59][16].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[59][16].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[59][16].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[59][16].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[59][16].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[59][16].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[59][16].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[59][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[59][16].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[59][17].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[59][17].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[59][17].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[59][17].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[59][17].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[59][17].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[59][17].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[59][17].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[59][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[59][17].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[59][18].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[59][18].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[59][18].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[59][18].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[59][18].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[59][18].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[59][18].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[59][18].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[59][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[59][18].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[59][19].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[59][19].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[59][19].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[59][19].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[59][19].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[59][19].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[59][19].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[59][19].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[59][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[59][19].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[59][20].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[59][20].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[59][20].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[59][20].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[59][20].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[59][20].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[59][20].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[59][20].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[59][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[59][20].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[59][21].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[59][21].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[59][21].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[59][21].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[59][21].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[59][21].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[59][21].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[59][21].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[59][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[59][21].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[59][22].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[59][22].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[59][22].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[59][22].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[59][22].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[59][22].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[59][22].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[59][22].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[59][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[59][22].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[59][23].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[59][23].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[59][23].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[59][23].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[59][23].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[59][23].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[59][23].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[59][23].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[59][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[59][23].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[59][24].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[59][24].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[59][24].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[59][24].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[59][24].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[59][24].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[59][24].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[59][24].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[59][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[59][24].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[59][25].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[59][25].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[59][25].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[59][25].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[59][25].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[59][25].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[59][25].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[59][25].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[59][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[59][25].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[59][26].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[59][26].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[59][26].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[59][26].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[59][26].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[59][26].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[59][26].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[59][26].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[59][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[59][26].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[59][27].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[59][27].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[59][27].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[59][27].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[59][27].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[59][27].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[59][27].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[59][27].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[59][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[59][27].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[59][28].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[59][28].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[59][28].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[59][28].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[59][28].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[59][28].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[59][28].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[59][28].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[59][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[59][28].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[59][29].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[59][29].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[59][29].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[59][29].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[59][29].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[59][29].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[59][29].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[59][29].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[59][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[59][29].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[59][30].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[59][30].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[59][30].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[59][30].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[59][30].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[59][30].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[59][30].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[59][30].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[59][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[59][30].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[59][31].dma__memc__write_valid      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[59][31].dma__memc__write_address    = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[59][31].dma__memc__write_data       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[59][31].dma__memc__read_valid       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[59][31].dma__memc__read_address     = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[59][31].dma__memc__read_pause       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[59][31].memc__dma__write_ready      = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[59][31].memc__dma__read_data        = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[59][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[59][31].memc__dma__read_ready       = pe_array_inst.pe_inst[59].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 60
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[60][0].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[60][0].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[60][0].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[60][0].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[60][0].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[60][0].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[60][0].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[60][0].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[60][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[60][0].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[60][1].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[60][1].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[60][1].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[60][1].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[60][1].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[60][1].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[60][1].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[60][1].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[60][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[60][1].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[60][2].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[60][2].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[60][2].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[60][2].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[60][2].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[60][2].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[60][2].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[60][2].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[60][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[60][2].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[60][3].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[60][3].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[60][3].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[60][3].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[60][3].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[60][3].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[60][3].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[60][3].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[60][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[60][3].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[60][4].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[60][4].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[60][4].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[60][4].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[60][4].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[60][4].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[60][4].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[60][4].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[60][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[60][4].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[60][5].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[60][5].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[60][5].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[60][5].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[60][5].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[60][5].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[60][5].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[60][5].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[60][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[60][5].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[60][6].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[60][6].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[60][6].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[60][6].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[60][6].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[60][6].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[60][6].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[60][6].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[60][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[60][6].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[60][7].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[60][7].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[60][7].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[60][7].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[60][7].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[60][7].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[60][7].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[60][7].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[60][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[60][7].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[60][8].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[60][8].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[60][8].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[60][8].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[60][8].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[60][8].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[60][8].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[60][8].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[60][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[60][8].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[60][9].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[60][9].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[60][9].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[60][9].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[60][9].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[60][9].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[60][9].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[60][9].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[60][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[60][9].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[60][10].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[60][10].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[60][10].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[60][10].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[60][10].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[60][10].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[60][10].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[60][10].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[60][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[60][10].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[60][11].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[60][11].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[60][11].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[60][11].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[60][11].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[60][11].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[60][11].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[60][11].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[60][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[60][11].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[60][12].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[60][12].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[60][12].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[60][12].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[60][12].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[60][12].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[60][12].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[60][12].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[60][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[60][12].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[60][13].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[60][13].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[60][13].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[60][13].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[60][13].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[60][13].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[60][13].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[60][13].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[60][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[60][13].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[60][14].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[60][14].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[60][14].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[60][14].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[60][14].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[60][14].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[60][14].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[60][14].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[60][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[60][14].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[60][15].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[60][15].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[60][15].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[60][15].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[60][15].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[60][15].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[60][15].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[60][15].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[60][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[60][15].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[60][16].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[60][16].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[60][16].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[60][16].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[60][16].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[60][16].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[60][16].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[60][16].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[60][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[60][16].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[60][17].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[60][17].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[60][17].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[60][17].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[60][17].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[60][17].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[60][17].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[60][17].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[60][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[60][17].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[60][18].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[60][18].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[60][18].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[60][18].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[60][18].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[60][18].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[60][18].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[60][18].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[60][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[60][18].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[60][19].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[60][19].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[60][19].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[60][19].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[60][19].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[60][19].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[60][19].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[60][19].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[60][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[60][19].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[60][20].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[60][20].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[60][20].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[60][20].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[60][20].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[60][20].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[60][20].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[60][20].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[60][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[60][20].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[60][21].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[60][21].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[60][21].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[60][21].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[60][21].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[60][21].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[60][21].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[60][21].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[60][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[60][21].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[60][22].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[60][22].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[60][22].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[60][22].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[60][22].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[60][22].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[60][22].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[60][22].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[60][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[60][22].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[60][23].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[60][23].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[60][23].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[60][23].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[60][23].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[60][23].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[60][23].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[60][23].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[60][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[60][23].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[60][24].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[60][24].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[60][24].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[60][24].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[60][24].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[60][24].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[60][24].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[60][24].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[60][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[60][24].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[60][25].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[60][25].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[60][25].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[60][25].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[60][25].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[60][25].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[60][25].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[60][25].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[60][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[60][25].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[60][26].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[60][26].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[60][26].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[60][26].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[60][26].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[60][26].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[60][26].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[60][26].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[60][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[60][26].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[60][27].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[60][27].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[60][27].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[60][27].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[60][27].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[60][27].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[60][27].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[60][27].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[60][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[60][27].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[60][28].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[60][28].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[60][28].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[60][28].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[60][28].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[60][28].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[60][28].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[60][28].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[60][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[60][28].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[60][29].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[60][29].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[60][29].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[60][29].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[60][29].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[60][29].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[60][29].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[60][29].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[60][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[60][29].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[60][30].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[60][30].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[60][30].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[60][30].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[60][30].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[60][30].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[60][30].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[60][30].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[60][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[60][30].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[60][31].dma__memc__write_valid      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[60][31].dma__memc__write_address    = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[60][31].dma__memc__write_data       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[60][31].dma__memc__read_valid       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[60][31].dma__memc__read_address     = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[60][31].dma__memc__read_pause       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[60][31].memc__dma__write_ready      = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[60][31].memc__dma__read_data        = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[60][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[60][31].memc__dma__read_ready       = pe_array_inst.pe_inst[60].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 61
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[61][0].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[61][0].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[61][0].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[61][0].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[61][0].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[61][0].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[61][0].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[61][0].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[61][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[61][0].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[61][1].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[61][1].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[61][1].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[61][1].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[61][1].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[61][1].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[61][1].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[61][1].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[61][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[61][1].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[61][2].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[61][2].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[61][2].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[61][2].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[61][2].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[61][2].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[61][2].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[61][2].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[61][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[61][2].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[61][3].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[61][3].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[61][3].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[61][3].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[61][3].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[61][3].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[61][3].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[61][3].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[61][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[61][3].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[61][4].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[61][4].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[61][4].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[61][4].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[61][4].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[61][4].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[61][4].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[61][4].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[61][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[61][4].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[61][5].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[61][5].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[61][5].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[61][5].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[61][5].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[61][5].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[61][5].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[61][5].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[61][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[61][5].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[61][6].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[61][6].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[61][6].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[61][6].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[61][6].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[61][6].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[61][6].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[61][6].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[61][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[61][6].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[61][7].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[61][7].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[61][7].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[61][7].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[61][7].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[61][7].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[61][7].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[61][7].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[61][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[61][7].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[61][8].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[61][8].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[61][8].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[61][8].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[61][8].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[61][8].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[61][8].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[61][8].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[61][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[61][8].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[61][9].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[61][9].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[61][9].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[61][9].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[61][9].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[61][9].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[61][9].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[61][9].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[61][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[61][9].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[61][10].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[61][10].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[61][10].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[61][10].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[61][10].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[61][10].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[61][10].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[61][10].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[61][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[61][10].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[61][11].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[61][11].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[61][11].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[61][11].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[61][11].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[61][11].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[61][11].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[61][11].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[61][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[61][11].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[61][12].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[61][12].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[61][12].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[61][12].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[61][12].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[61][12].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[61][12].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[61][12].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[61][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[61][12].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[61][13].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[61][13].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[61][13].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[61][13].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[61][13].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[61][13].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[61][13].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[61][13].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[61][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[61][13].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[61][14].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[61][14].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[61][14].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[61][14].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[61][14].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[61][14].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[61][14].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[61][14].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[61][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[61][14].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[61][15].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[61][15].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[61][15].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[61][15].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[61][15].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[61][15].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[61][15].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[61][15].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[61][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[61][15].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[61][16].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[61][16].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[61][16].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[61][16].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[61][16].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[61][16].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[61][16].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[61][16].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[61][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[61][16].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[61][17].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[61][17].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[61][17].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[61][17].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[61][17].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[61][17].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[61][17].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[61][17].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[61][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[61][17].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[61][18].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[61][18].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[61][18].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[61][18].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[61][18].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[61][18].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[61][18].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[61][18].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[61][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[61][18].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[61][19].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[61][19].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[61][19].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[61][19].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[61][19].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[61][19].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[61][19].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[61][19].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[61][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[61][19].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[61][20].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[61][20].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[61][20].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[61][20].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[61][20].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[61][20].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[61][20].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[61][20].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[61][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[61][20].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[61][21].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[61][21].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[61][21].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[61][21].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[61][21].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[61][21].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[61][21].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[61][21].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[61][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[61][21].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[61][22].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[61][22].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[61][22].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[61][22].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[61][22].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[61][22].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[61][22].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[61][22].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[61][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[61][22].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[61][23].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[61][23].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[61][23].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[61][23].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[61][23].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[61][23].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[61][23].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[61][23].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[61][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[61][23].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[61][24].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[61][24].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[61][24].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[61][24].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[61][24].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[61][24].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[61][24].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[61][24].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[61][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[61][24].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[61][25].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[61][25].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[61][25].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[61][25].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[61][25].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[61][25].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[61][25].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[61][25].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[61][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[61][25].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[61][26].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[61][26].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[61][26].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[61][26].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[61][26].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[61][26].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[61][26].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[61][26].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[61][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[61][26].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[61][27].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[61][27].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[61][27].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[61][27].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[61][27].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[61][27].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[61][27].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[61][27].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[61][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[61][27].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[61][28].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[61][28].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[61][28].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[61][28].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[61][28].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[61][28].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[61][28].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[61][28].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[61][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[61][28].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[61][29].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[61][29].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[61][29].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[61][29].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[61][29].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[61][29].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[61][29].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[61][29].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[61][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[61][29].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[61][30].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[61][30].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[61][30].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[61][30].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[61][30].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[61][30].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[61][30].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[61][30].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[61][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[61][30].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[61][31].dma__memc__write_valid      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[61][31].dma__memc__write_address    = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[61][31].dma__memc__write_data       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[61][31].dma__memc__read_valid       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[61][31].dma__memc__read_address     = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[61][31].dma__memc__read_pause       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[61][31].memc__dma__write_ready      = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[61][31].memc__dma__read_data        = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[61][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[61][31].memc__dma__read_ready       = pe_array_inst.pe_inst[61].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 62
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[62][0].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[62][0].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[62][0].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[62][0].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[62][0].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[62][0].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[62][0].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[62][0].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[62][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[62][0].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[62][1].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[62][1].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[62][1].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[62][1].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[62][1].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[62][1].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[62][1].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[62][1].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[62][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[62][1].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[62][2].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[62][2].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[62][2].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[62][2].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[62][2].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[62][2].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[62][2].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[62][2].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[62][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[62][2].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[62][3].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[62][3].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[62][3].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[62][3].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[62][3].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[62][3].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[62][3].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[62][3].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[62][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[62][3].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[62][4].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[62][4].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[62][4].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[62][4].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[62][4].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[62][4].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[62][4].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[62][4].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[62][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[62][4].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[62][5].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[62][5].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[62][5].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[62][5].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[62][5].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[62][5].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[62][5].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[62][5].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[62][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[62][5].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[62][6].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[62][6].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[62][6].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[62][6].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[62][6].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[62][6].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[62][6].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[62][6].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[62][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[62][6].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[62][7].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[62][7].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[62][7].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[62][7].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[62][7].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[62][7].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[62][7].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[62][7].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[62][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[62][7].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[62][8].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[62][8].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[62][8].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[62][8].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[62][8].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[62][8].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[62][8].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[62][8].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[62][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[62][8].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[62][9].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[62][9].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[62][9].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[62][9].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[62][9].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[62][9].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[62][9].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[62][9].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[62][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[62][9].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[62][10].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[62][10].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[62][10].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[62][10].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[62][10].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[62][10].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[62][10].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[62][10].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[62][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[62][10].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[62][11].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[62][11].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[62][11].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[62][11].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[62][11].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[62][11].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[62][11].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[62][11].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[62][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[62][11].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[62][12].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[62][12].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[62][12].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[62][12].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[62][12].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[62][12].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[62][12].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[62][12].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[62][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[62][12].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[62][13].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[62][13].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[62][13].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[62][13].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[62][13].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[62][13].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[62][13].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[62][13].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[62][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[62][13].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[62][14].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[62][14].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[62][14].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[62][14].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[62][14].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[62][14].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[62][14].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[62][14].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[62][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[62][14].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[62][15].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[62][15].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[62][15].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[62][15].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[62][15].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[62][15].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[62][15].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[62][15].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[62][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[62][15].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[62][16].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[62][16].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[62][16].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[62][16].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[62][16].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[62][16].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[62][16].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[62][16].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[62][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[62][16].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[62][17].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[62][17].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[62][17].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[62][17].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[62][17].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[62][17].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[62][17].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[62][17].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[62][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[62][17].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[62][18].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[62][18].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[62][18].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[62][18].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[62][18].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[62][18].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[62][18].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[62][18].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[62][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[62][18].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[62][19].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[62][19].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[62][19].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[62][19].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[62][19].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[62][19].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[62][19].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[62][19].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[62][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[62][19].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[62][20].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[62][20].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[62][20].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[62][20].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[62][20].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[62][20].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[62][20].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[62][20].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[62][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[62][20].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[62][21].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[62][21].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[62][21].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[62][21].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[62][21].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[62][21].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[62][21].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[62][21].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[62][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[62][21].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[62][22].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[62][22].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[62][22].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[62][22].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[62][22].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[62][22].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[62][22].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[62][22].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[62][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[62][22].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[62][23].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[62][23].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[62][23].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[62][23].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[62][23].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[62][23].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[62][23].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[62][23].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[62][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[62][23].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[62][24].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[62][24].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[62][24].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[62][24].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[62][24].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[62][24].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[62][24].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[62][24].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[62][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[62][24].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[62][25].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[62][25].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[62][25].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[62][25].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[62][25].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[62][25].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[62][25].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[62][25].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[62][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[62][25].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[62][26].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[62][26].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[62][26].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[62][26].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[62][26].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[62][26].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[62][26].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[62][26].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[62][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[62][26].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[62][27].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[62][27].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[62][27].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[62][27].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[62][27].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[62][27].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[62][27].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[62][27].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[62][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[62][27].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[62][28].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[62][28].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[62][28].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[62][28].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[62][28].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[62][28].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[62][28].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[62][28].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[62][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[62][28].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[62][29].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[62][29].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[62][29].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[62][29].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[62][29].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[62][29].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[62][29].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[62][29].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[62][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[62][29].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[62][30].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[62][30].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[62][30].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[62][30].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[62][30].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[62][30].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[62][30].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[62][30].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[62][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[62][30].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[62][31].dma__memc__write_valid      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[62][31].dma__memc__write_address    = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[62][31].dma__memc__write_data       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[62][31].dma__memc__read_valid       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[62][31].dma__memc__read_address     = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[62][31].dma__memc__read_pause       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[62][31].memc__dma__write_ready      = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[62][31].memc__dma__read_data        = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[62][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[62][31].memc__dma__read_ready       = pe_array_inst.pe_inst[62].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 63
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[63][0].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[63][0].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[63][0].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[63][0].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[63][0].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[63][0].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[63][0].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[63][0].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[63][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[63][0].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[63][1].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[63][1].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[63][1].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[63][1].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[63][1].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[63][1].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[63][1].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[63][1].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[63][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[63][1].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[63][2].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[63][2].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[63][2].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[63][2].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[63][2].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[63][2].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[63][2].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[63][2].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[63][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[63][2].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[63][3].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[63][3].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[63][3].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[63][3].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[63][3].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[63][3].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[63][3].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[63][3].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[63][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[63][3].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[63][4].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[63][4].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[63][4].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[63][4].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[63][4].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[63][4].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[63][4].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[63][4].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[63][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[63][4].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[63][5].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[63][5].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[63][5].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[63][5].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[63][5].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[63][5].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[63][5].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[63][5].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[63][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[63][5].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[63][6].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[63][6].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[63][6].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[63][6].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[63][6].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[63][6].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[63][6].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[63][6].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[63][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[63][6].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[63][7].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[63][7].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[63][7].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[63][7].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[63][7].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[63][7].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[63][7].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[63][7].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[63][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[63][7].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[63][8].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[63][8].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[63][8].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[63][8].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[63][8].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[63][8].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[63][8].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[63][8].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[63][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[63][8].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[63][9].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[63][9].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[63][9].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[63][9].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[63][9].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[63][9].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[63][9].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[63][9].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[63][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[63][9].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[63][10].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[63][10].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[63][10].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[63][10].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[63][10].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[63][10].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[63][10].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[63][10].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[63][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[63][10].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[63][11].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[63][11].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[63][11].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[63][11].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[63][11].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[63][11].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[63][11].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[63][11].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[63][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[63][11].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[63][12].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[63][12].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[63][12].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[63][12].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[63][12].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[63][12].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[63][12].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[63][12].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[63][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[63][12].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[63][13].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[63][13].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[63][13].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[63][13].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[63][13].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[63][13].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[63][13].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[63][13].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[63][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[63][13].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[63][14].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[63][14].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[63][14].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[63][14].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[63][14].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[63][14].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[63][14].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[63][14].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[63][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[63][14].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[63][15].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[63][15].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[63][15].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[63][15].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[63][15].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[63][15].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[63][15].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[63][15].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[63][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[63][15].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[63][16].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[63][16].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[63][16].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[63][16].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[63][16].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[63][16].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[63][16].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[63][16].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[63][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[63][16].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[63][17].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[63][17].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[63][17].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[63][17].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[63][17].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[63][17].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[63][17].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[63][17].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[63][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[63][17].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[63][18].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[63][18].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[63][18].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[63][18].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[63][18].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[63][18].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[63][18].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[63][18].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[63][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[63][18].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[63][19].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[63][19].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[63][19].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[63][19].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[63][19].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[63][19].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[63][19].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[63][19].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[63][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[63][19].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[63][20].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[63][20].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[63][20].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[63][20].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[63][20].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[63][20].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[63][20].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[63][20].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[63][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[63][20].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[63][21].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[63][21].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[63][21].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[63][21].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[63][21].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[63][21].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[63][21].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[63][21].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[63][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[63][21].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[63][22].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[63][22].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[63][22].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[63][22].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[63][22].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[63][22].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[63][22].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[63][22].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[63][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[63][22].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[63][23].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[63][23].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[63][23].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[63][23].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[63][23].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[63][23].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[63][23].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[63][23].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[63][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[63][23].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[63][24].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[63][24].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[63][24].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[63][24].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[63][24].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[63][24].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[63][24].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[63][24].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[63][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[63][24].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[63][25].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[63][25].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[63][25].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[63][25].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[63][25].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[63][25].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[63][25].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[63][25].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[63][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[63][25].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[63][26].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[63][26].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[63][26].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[63][26].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[63][26].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[63][26].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[63][26].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[63][26].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[63][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[63][26].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[63][27].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[63][27].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[63][27].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[63][27].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[63][27].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[63][27].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[63][27].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[63][27].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[63][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[63][27].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[63][28].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[63][28].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[63][28].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[63][28].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[63][28].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[63][28].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[63][28].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[63][28].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[63][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[63][28].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[63][29].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[63][29].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[63][29].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[63][29].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[63][29].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[63][29].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[63][29].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[63][29].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[63][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[63][29].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[63][30].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[63][30].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[63][30].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[63][30].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[63][30].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[63][30].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[63][30].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[63][30].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[63][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[63][30].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[63][31].dma__memc__write_valid      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[63][31].dma__memc__write_address    = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[63][31].dma__memc__write_data       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[63][31].dma__memc__read_valid       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[63][31].dma__memc__read_address     = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[63][31].dma__memc__read_pause       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[63][31].memc__dma__write_ready      = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[63][31].memc__dma__read_data        = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[63][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[63][31].memc__dma__read_ready       = pe_array_inst.pe_inst[63].pe.mem_acc_cont.memc__dma__read_ready31         ;
