
  assign stOp_lane[0].reg__stOp__ready = reg__sdp__lane0_ready          ;
  assign sdp__reg__lane0_valid         = stOp_lane[0].stOp__reg__valid  ;
  assign sdp__reg__lane0_data          = stOp_lane[0].stOp__reg__data   ;
  assign stOp_lane[1].reg__stOp__ready = reg__sdp__lane1_ready          ;
  assign sdp__reg__lane1_valid         = stOp_lane[1].stOp__reg__valid  ;
  assign sdp__reg__lane1_data          = stOp_lane[1].stOp__reg__data   ;
  assign stOp_lane[2].reg__stOp__ready = reg__sdp__lane2_ready          ;
  assign sdp__reg__lane2_valid         = stOp_lane[2].stOp__reg__valid  ;
  assign sdp__reg__lane2_data          = stOp_lane[2].stOp__reg__data   ;
  assign stOp_lane[3].reg__stOp__ready = reg__sdp__lane3_ready          ;
  assign sdp__reg__lane3_valid         = stOp_lane[3].stOp__reg__valid  ;
  assign sdp__reg__lane3_data          = stOp_lane[3].stOp__reg__data   ;
  assign stOp_lane[4].reg__stOp__ready = reg__sdp__lane4_ready          ;
  assign sdp__reg__lane4_valid         = stOp_lane[4].stOp__reg__valid  ;
  assign sdp__reg__lane4_data          = stOp_lane[4].stOp__reg__data   ;
  assign stOp_lane[5].reg__stOp__ready = reg__sdp__lane5_ready          ;
  assign sdp__reg__lane5_valid         = stOp_lane[5].stOp__reg__valid  ;
  assign sdp__reg__lane5_data          = stOp_lane[5].stOp__reg__data   ;
  assign stOp_lane[6].reg__stOp__ready = reg__sdp__lane6_ready          ;
  assign sdp__reg__lane6_valid         = stOp_lane[6].stOp__reg__valid  ;
  assign sdp__reg__lane6_data          = stOp_lane[6].stOp__reg__data   ;
  assign stOp_lane[7].reg__stOp__ready = reg__sdp__lane7_ready          ;
  assign sdp__reg__lane7_valid         = stOp_lane[7].stOp__reg__valid  ;
  assign sdp__reg__lane7_data          = stOp_lane[7].stOp__reg__data   ;
  assign stOp_lane[8].reg__stOp__ready = reg__sdp__lane8_ready          ;
  assign sdp__reg__lane8_valid         = stOp_lane[8].stOp__reg__valid  ;
  assign sdp__reg__lane8_data          = stOp_lane[8].stOp__reg__data   ;
  assign stOp_lane[9].reg__stOp__ready = reg__sdp__lane9_ready          ;
  assign sdp__reg__lane9_valid         = stOp_lane[9].stOp__reg__valid  ;
  assign sdp__reg__lane9_data          = stOp_lane[9].stOp__reg__data   ;
  assign stOp_lane[10].reg__stOp__ready = reg__sdp__lane10_ready          ;
  assign sdp__reg__lane10_valid         = stOp_lane[10].stOp__reg__valid  ;
  assign sdp__reg__lane10_data          = stOp_lane[10].stOp__reg__data   ;
  assign stOp_lane[11].reg__stOp__ready = reg__sdp__lane11_ready          ;
  assign sdp__reg__lane11_valid         = stOp_lane[11].stOp__reg__valid  ;
  assign sdp__reg__lane11_data          = stOp_lane[11].stOp__reg__data   ;
  assign stOp_lane[12].reg__stOp__ready = reg__sdp__lane12_ready          ;
  assign sdp__reg__lane12_valid         = stOp_lane[12].stOp__reg__valid  ;
  assign sdp__reg__lane12_data          = stOp_lane[12].stOp__reg__data   ;
  assign stOp_lane[13].reg__stOp__ready = reg__sdp__lane13_ready          ;
  assign sdp__reg__lane13_valid         = stOp_lane[13].stOp__reg__valid  ;
  assign sdp__reg__lane13_data          = stOp_lane[13].stOp__reg__data   ;
  assign stOp_lane[14].reg__stOp__ready = reg__sdp__lane14_ready          ;
  assign sdp__reg__lane14_valid         = stOp_lane[14].stOp__reg__valid  ;
  assign sdp__reg__lane14_data          = stOp_lane[14].stOp__reg__data   ;
  assign stOp_lane[15].reg__stOp__ready = reg__sdp__lane15_ready          ;
  assign sdp__reg__lane15_valid         = stOp_lane[15].stOp__reg__valid  ;
  assign sdp__reg__lane15_data          = stOp_lane[15].stOp__reg__data   ;
  assign stOp_lane[16].reg__stOp__ready = reg__sdp__lane16_ready          ;
  assign sdp__reg__lane16_valid         = stOp_lane[16].stOp__reg__valid  ;
  assign sdp__reg__lane16_data          = stOp_lane[16].stOp__reg__data   ;
  assign stOp_lane[17].reg__stOp__ready = reg__sdp__lane17_ready          ;
  assign sdp__reg__lane17_valid         = stOp_lane[17].stOp__reg__valid  ;
  assign sdp__reg__lane17_data          = stOp_lane[17].stOp__reg__data   ;
  assign stOp_lane[18].reg__stOp__ready = reg__sdp__lane18_ready          ;
  assign sdp__reg__lane18_valid         = stOp_lane[18].stOp__reg__valid  ;
  assign sdp__reg__lane18_data          = stOp_lane[18].stOp__reg__data   ;
  assign stOp_lane[19].reg__stOp__ready = reg__sdp__lane19_ready          ;
  assign sdp__reg__lane19_valid         = stOp_lane[19].stOp__reg__valid  ;
  assign sdp__reg__lane19_data          = stOp_lane[19].stOp__reg__data   ;
  assign stOp_lane[20].reg__stOp__ready = reg__sdp__lane20_ready          ;
  assign sdp__reg__lane20_valid         = stOp_lane[20].stOp__reg__valid  ;
  assign sdp__reg__lane20_data          = stOp_lane[20].stOp__reg__data   ;
  assign stOp_lane[21].reg__stOp__ready = reg__sdp__lane21_ready          ;
  assign sdp__reg__lane21_valid         = stOp_lane[21].stOp__reg__valid  ;
  assign sdp__reg__lane21_data          = stOp_lane[21].stOp__reg__data   ;
  assign stOp_lane[22].reg__stOp__ready = reg__sdp__lane22_ready          ;
  assign sdp__reg__lane22_valid         = stOp_lane[22].stOp__reg__valid  ;
  assign sdp__reg__lane22_data          = stOp_lane[22].stOp__reg__data   ;
  assign stOp_lane[23].reg__stOp__ready = reg__sdp__lane23_ready          ;
  assign sdp__reg__lane23_valid         = stOp_lane[23].stOp__reg__valid  ;
  assign sdp__reg__lane23_data          = stOp_lane[23].stOp__reg__data   ;
  assign stOp_lane[24].reg__stOp__ready = reg__sdp__lane24_ready          ;
  assign sdp__reg__lane24_valid         = stOp_lane[24].stOp__reg__valid  ;
  assign sdp__reg__lane24_data          = stOp_lane[24].stOp__reg__data   ;
  assign stOp_lane[25].reg__stOp__ready = reg__sdp__lane25_ready          ;
  assign sdp__reg__lane25_valid         = stOp_lane[25].stOp__reg__valid  ;
  assign sdp__reg__lane25_data          = stOp_lane[25].stOp__reg__data   ;
  assign stOp_lane[26].reg__stOp__ready = reg__sdp__lane26_ready          ;
  assign sdp__reg__lane26_valid         = stOp_lane[26].stOp__reg__valid  ;
  assign sdp__reg__lane26_data          = stOp_lane[26].stOp__reg__data   ;
  assign stOp_lane[27].reg__stOp__ready = reg__sdp__lane27_ready          ;
  assign sdp__reg__lane27_valid         = stOp_lane[27].stOp__reg__valid  ;
  assign sdp__reg__lane27_data          = stOp_lane[27].stOp__reg__data   ;
  assign stOp_lane[28].reg__stOp__ready = reg__sdp__lane28_ready          ;
  assign sdp__reg__lane28_valid         = stOp_lane[28].stOp__reg__valid  ;
  assign sdp__reg__lane28_data          = stOp_lane[28].stOp__reg__data   ;
  assign stOp_lane[29].reg__stOp__ready = reg__sdp__lane29_ready          ;
  assign sdp__reg__lane29_valid         = stOp_lane[29].stOp__reg__valid  ;
  assign sdp__reg__lane29_data          = stOp_lane[29].stOp__reg__data   ;
  assign stOp_lane[30].reg__stOp__ready = reg__sdp__lane30_ready          ;
  assign sdp__reg__lane30_valid         = stOp_lane[30].stOp__reg__valid  ;
  assign sdp__reg__lane30_data          = stOp_lane[30].stOp__reg__data   ;
  assign stOp_lane[31].reg__stOp__ready = reg__sdp__lane31_ready          ;
  assign sdp__reg__lane31_valid         = stOp_lane[31].stOp__reg__valid  ;
  assign sdp__reg__lane31_data          = stOp_lane[31].stOp__reg__data   ;

  assign reg__sdp__lane0_ready  = 1'b1          ;
  assign reg__sdp__lane1_ready  = 1'b1          ;
  assign reg__sdp__lane2_ready  = 1'b1          ;
  assign reg__sdp__lane3_ready  = 1'b1          ;
  assign reg__sdp__lane4_ready  = 1'b1          ;
  assign reg__sdp__lane5_ready  = 1'b1          ;
  assign reg__sdp__lane6_ready  = 1'b1          ;
  assign reg__sdp__lane7_ready  = 1'b1          ;
  assign reg__sdp__lane8_ready  = 1'b1          ;
  assign reg__sdp__lane9_ready  = 1'b1          ;
  assign reg__sdp__lane10_ready  = 1'b1          ;
  assign reg__sdp__lane11_ready  = 1'b1          ;
  assign reg__sdp__lane12_ready  = 1'b1          ;
  assign reg__sdp__lane13_ready  = 1'b1          ;
  assign reg__sdp__lane14_ready  = 1'b1          ;
  assign reg__sdp__lane15_ready  = 1'b1          ;
  assign reg__sdp__lane16_ready  = 1'b1          ;
  assign reg__sdp__lane17_ready  = 1'b1          ;
  assign reg__sdp__lane18_ready  = 1'b1          ;
  assign reg__sdp__lane19_ready  = 1'b1          ;
  assign reg__sdp__lane20_ready  = 1'b1          ;
  assign reg__sdp__lane21_ready  = 1'b1          ;
  assign reg__sdp__lane22_ready  = 1'b1          ;
  assign reg__sdp__lane23_ready  = 1'b1          ;
  assign reg__sdp__lane24_ready  = 1'b1          ;
  assign reg__sdp__lane25_ready  = 1'b1          ;
  assign reg__sdp__lane26_ready  = 1'b1          ;
  assign reg__sdp__lane27_ready  = 1'b1          ;
  assign reg__sdp__lane28_ready  = 1'b1          ;
  assign reg__sdp__lane29_ready  = 1'b1          ;
  assign reg__sdp__lane30_ready  = 1'b1          ;
  assign reg__sdp__lane31_ready  = 1'b1          ;
