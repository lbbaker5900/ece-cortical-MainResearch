
  input                                         std__mgr0__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane0_strm0_data        ;
  output                                        mgr0__std__lane0_strm0_data_valid  ;

  input                                         std__mgr0__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane0_strm1_data        ;
  output                                        mgr0__std__lane0_strm1_data_valid  ;

  input                                         std__mgr0__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane1_strm0_data        ;
  output                                        mgr0__std__lane1_strm0_data_valid  ;

  input                                         std__mgr0__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane1_strm1_data        ;
  output                                        mgr0__std__lane1_strm1_data_valid  ;

  input                                         std__mgr0__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane2_strm0_data        ;
  output                                        mgr0__std__lane2_strm0_data_valid  ;

  input                                         std__mgr0__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane2_strm1_data        ;
  output                                        mgr0__std__lane2_strm1_data_valid  ;

  input                                         std__mgr0__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane3_strm0_data        ;
  output                                        mgr0__std__lane3_strm0_data_valid  ;

  input                                         std__mgr0__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane3_strm1_data        ;
  output                                        mgr0__std__lane3_strm1_data_valid  ;

  input                                         std__mgr0__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane4_strm0_data        ;
  output                                        mgr0__std__lane4_strm0_data_valid  ;

  input                                         std__mgr0__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane4_strm1_data        ;
  output                                        mgr0__std__lane4_strm1_data_valid  ;

  input                                         std__mgr0__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane5_strm0_data        ;
  output                                        mgr0__std__lane5_strm0_data_valid  ;

  input                                         std__mgr0__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane5_strm1_data        ;
  output                                        mgr0__std__lane5_strm1_data_valid  ;

  input                                         std__mgr0__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane6_strm0_data        ;
  output                                        mgr0__std__lane6_strm0_data_valid  ;

  input                                         std__mgr0__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane6_strm1_data        ;
  output                                        mgr0__std__lane6_strm1_data_valid  ;

  input                                         std__mgr0__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane7_strm0_data        ;
  output                                        mgr0__std__lane7_strm0_data_valid  ;

  input                                         std__mgr0__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane7_strm1_data        ;
  output                                        mgr0__std__lane7_strm1_data_valid  ;

  input                                         std__mgr0__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane8_strm0_data        ;
  output                                        mgr0__std__lane8_strm0_data_valid  ;

  input                                         std__mgr0__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane8_strm1_data        ;
  output                                        mgr0__std__lane8_strm1_data_valid  ;

  input                                         std__mgr0__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane9_strm0_data        ;
  output                                        mgr0__std__lane9_strm0_data_valid  ;

  input                                         std__mgr0__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane9_strm1_data        ;
  output                                        mgr0__std__lane9_strm1_data_valid  ;

  input                                         std__mgr0__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane10_strm0_data        ;
  output                                        mgr0__std__lane10_strm0_data_valid  ;

  input                                         std__mgr0__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane10_strm1_data        ;
  output                                        mgr0__std__lane10_strm1_data_valid  ;

  input                                         std__mgr0__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane11_strm0_data        ;
  output                                        mgr0__std__lane11_strm0_data_valid  ;

  input                                         std__mgr0__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane11_strm1_data        ;
  output                                        mgr0__std__lane11_strm1_data_valid  ;

  input                                         std__mgr0__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane12_strm0_data        ;
  output                                        mgr0__std__lane12_strm0_data_valid  ;

  input                                         std__mgr0__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane12_strm1_data        ;
  output                                        mgr0__std__lane12_strm1_data_valid  ;

  input                                         std__mgr0__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane13_strm0_data        ;
  output                                        mgr0__std__lane13_strm0_data_valid  ;

  input                                         std__mgr0__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane13_strm1_data        ;
  output                                        mgr0__std__lane13_strm1_data_valid  ;

  input                                         std__mgr0__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane14_strm0_data        ;
  output                                        mgr0__std__lane14_strm0_data_valid  ;

  input                                         std__mgr0__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane14_strm1_data        ;
  output                                        mgr0__std__lane14_strm1_data_valid  ;

  input                                         std__mgr0__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane15_strm0_data        ;
  output                                        mgr0__std__lane15_strm0_data_valid  ;

  input                                         std__mgr0__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane15_strm1_data        ;
  output                                        mgr0__std__lane15_strm1_data_valid  ;

  input                                         std__mgr0__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane16_strm0_data        ;
  output                                        mgr0__std__lane16_strm0_data_valid  ;

  input                                         std__mgr0__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane16_strm1_data        ;
  output                                        mgr0__std__lane16_strm1_data_valid  ;

  input                                         std__mgr0__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane17_strm0_data        ;
  output                                        mgr0__std__lane17_strm0_data_valid  ;

  input                                         std__mgr0__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane17_strm1_data        ;
  output                                        mgr0__std__lane17_strm1_data_valid  ;

  input                                         std__mgr0__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane18_strm0_data        ;
  output                                        mgr0__std__lane18_strm0_data_valid  ;

  input                                         std__mgr0__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane18_strm1_data        ;
  output                                        mgr0__std__lane18_strm1_data_valid  ;

  input                                         std__mgr0__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane19_strm0_data        ;
  output                                        mgr0__std__lane19_strm0_data_valid  ;

  input                                         std__mgr0__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane19_strm1_data        ;
  output                                        mgr0__std__lane19_strm1_data_valid  ;

  input                                         std__mgr0__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane20_strm0_data        ;
  output                                        mgr0__std__lane20_strm0_data_valid  ;

  input                                         std__mgr0__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane20_strm1_data        ;
  output                                        mgr0__std__lane20_strm1_data_valid  ;

  input                                         std__mgr0__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane21_strm0_data        ;
  output                                        mgr0__std__lane21_strm0_data_valid  ;

  input                                         std__mgr0__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane21_strm1_data        ;
  output                                        mgr0__std__lane21_strm1_data_valid  ;

  input                                         std__mgr0__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane22_strm0_data        ;
  output                                        mgr0__std__lane22_strm0_data_valid  ;

  input                                         std__mgr0__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane22_strm1_data        ;
  output                                        mgr0__std__lane22_strm1_data_valid  ;

  input                                         std__mgr0__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane23_strm0_data        ;
  output                                        mgr0__std__lane23_strm0_data_valid  ;

  input                                         std__mgr0__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane23_strm1_data        ;
  output                                        mgr0__std__lane23_strm1_data_valid  ;

  input                                         std__mgr0__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane24_strm0_data        ;
  output                                        mgr0__std__lane24_strm0_data_valid  ;

  input                                         std__mgr0__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane24_strm1_data        ;
  output                                        mgr0__std__lane24_strm1_data_valid  ;

  input                                         std__mgr0__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane25_strm0_data        ;
  output                                        mgr0__std__lane25_strm0_data_valid  ;

  input                                         std__mgr0__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane25_strm1_data        ;
  output                                        mgr0__std__lane25_strm1_data_valid  ;

  input                                         std__mgr0__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane26_strm0_data        ;
  output                                        mgr0__std__lane26_strm0_data_valid  ;

  input                                         std__mgr0__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane26_strm1_data        ;
  output                                        mgr0__std__lane26_strm1_data_valid  ;

  input                                         std__mgr0__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane27_strm0_data        ;
  output                                        mgr0__std__lane27_strm0_data_valid  ;

  input                                         std__mgr0__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane27_strm1_data        ;
  output                                        mgr0__std__lane27_strm1_data_valid  ;

  input                                         std__mgr0__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane28_strm0_data        ;
  output                                        mgr0__std__lane28_strm0_data_valid  ;

  input                                         std__mgr0__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane28_strm1_data        ;
  output                                        mgr0__std__lane28_strm1_data_valid  ;

  input                                         std__mgr0__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane29_strm0_data        ;
  output                                        mgr0__std__lane29_strm0_data_valid  ;

  input                                         std__mgr0__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane29_strm1_data        ;
  output                                        mgr0__std__lane29_strm1_data_valid  ;

  input                                         std__mgr0__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane30_strm0_data        ;
  output                                        mgr0__std__lane30_strm0_data_valid  ;

  input                                         std__mgr0__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane30_strm1_data        ;
  output                                        mgr0__std__lane30_strm1_data_valid  ;

  input                                         std__mgr0__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane31_strm0_data        ;
  output                                        mgr0__std__lane31_strm0_data_valid  ;

  input                                         std__mgr0__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane31_strm1_data        ;
  output                                        mgr0__std__lane31_strm1_data_valid  ;

  input                                         std__mgr1__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane0_strm0_data        ;
  output                                        mgr1__std__lane0_strm0_data_valid  ;

  input                                         std__mgr1__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane0_strm1_data        ;
  output                                        mgr1__std__lane0_strm1_data_valid  ;

  input                                         std__mgr1__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane1_strm0_data        ;
  output                                        mgr1__std__lane1_strm0_data_valid  ;

  input                                         std__mgr1__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane1_strm1_data        ;
  output                                        mgr1__std__lane1_strm1_data_valid  ;

  input                                         std__mgr1__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane2_strm0_data        ;
  output                                        mgr1__std__lane2_strm0_data_valid  ;

  input                                         std__mgr1__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane2_strm1_data        ;
  output                                        mgr1__std__lane2_strm1_data_valid  ;

  input                                         std__mgr1__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane3_strm0_data        ;
  output                                        mgr1__std__lane3_strm0_data_valid  ;

  input                                         std__mgr1__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane3_strm1_data        ;
  output                                        mgr1__std__lane3_strm1_data_valid  ;

  input                                         std__mgr1__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane4_strm0_data        ;
  output                                        mgr1__std__lane4_strm0_data_valid  ;

  input                                         std__mgr1__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane4_strm1_data        ;
  output                                        mgr1__std__lane4_strm1_data_valid  ;

  input                                         std__mgr1__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane5_strm0_data        ;
  output                                        mgr1__std__lane5_strm0_data_valid  ;

  input                                         std__mgr1__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane5_strm1_data        ;
  output                                        mgr1__std__lane5_strm1_data_valid  ;

  input                                         std__mgr1__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane6_strm0_data        ;
  output                                        mgr1__std__lane6_strm0_data_valid  ;

  input                                         std__mgr1__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane6_strm1_data        ;
  output                                        mgr1__std__lane6_strm1_data_valid  ;

  input                                         std__mgr1__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane7_strm0_data        ;
  output                                        mgr1__std__lane7_strm0_data_valid  ;

  input                                         std__mgr1__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane7_strm1_data        ;
  output                                        mgr1__std__lane7_strm1_data_valid  ;

  input                                         std__mgr1__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane8_strm0_data        ;
  output                                        mgr1__std__lane8_strm0_data_valid  ;

  input                                         std__mgr1__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane8_strm1_data        ;
  output                                        mgr1__std__lane8_strm1_data_valid  ;

  input                                         std__mgr1__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane9_strm0_data        ;
  output                                        mgr1__std__lane9_strm0_data_valid  ;

  input                                         std__mgr1__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane9_strm1_data        ;
  output                                        mgr1__std__lane9_strm1_data_valid  ;

  input                                         std__mgr1__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane10_strm0_data        ;
  output                                        mgr1__std__lane10_strm0_data_valid  ;

  input                                         std__mgr1__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane10_strm1_data        ;
  output                                        mgr1__std__lane10_strm1_data_valid  ;

  input                                         std__mgr1__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane11_strm0_data        ;
  output                                        mgr1__std__lane11_strm0_data_valid  ;

  input                                         std__mgr1__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane11_strm1_data        ;
  output                                        mgr1__std__lane11_strm1_data_valid  ;

  input                                         std__mgr1__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane12_strm0_data        ;
  output                                        mgr1__std__lane12_strm0_data_valid  ;

  input                                         std__mgr1__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane12_strm1_data        ;
  output                                        mgr1__std__lane12_strm1_data_valid  ;

  input                                         std__mgr1__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane13_strm0_data        ;
  output                                        mgr1__std__lane13_strm0_data_valid  ;

  input                                         std__mgr1__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane13_strm1_data        ;
  output                                        mgr1__std__lane13_strm1_data_valid  ;

  input                                         std__mgr1__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane14_strm0_data        ;
  output                                        mgr1__std__lane14_strm0_data_valid  ;

  input                                         std__mgr1__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane14_strm1_data        ;
  output                                        mgr1__std__lane14_strm1_data_valid  ;

  input                                         std__mgr1__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane15_strm0_data        ;
  output                                        mgr1__std__lane15_strm0_data_valid  ;

  input                                         std__mgr1__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane15_strm1_data        ;
  output                                        mgr1__std__lane15_strm1_data_valid  ;

  input                                         std__mgr1__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane16_strm0_data        ;
  output                                        mgr1__std__lane16_strm0_data_valid  ;

  input                                         std__mgr1__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane16_strm1_data        ;
  output                                        mgr1__std__lane16_strm1_data_valid  ;

  input                                         std__mgr1__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane17_strm0_data        ;
  output                                        mgr1__std__lane17_strm0_data_valid  ;

  input                                         std__mgr1__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane17_strm1_data        ;
  output                                        mgr1__std__lane17_strm1_data_valid  ;

  input                                         std__mgr1__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane18_strm0_data        ;
  output                                        mgr1__std__lane18_strm0_data_valid  ;

  input                                         std__mgr1__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane18_strm1_data        ;
  output                                        mgr1__std__lane18_strm1_data_valid  ;

  input                                         std__mgr1__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane19_strm0_data        ;
  output                                        mgr1__std__lane19_strm0_data_valid  ;

  input                                         std__mgr1__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane19_strm1_data        ;
  output                                        mgr1__std__lane19_strm1_data_valid  ;

  input                                         std__mgr1__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane20_strm0_data        ;
  output                                        mgr1__std__lane20_strm0_data_valid  ;

  input                                         std__mgr1__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane20_strm1_data        ;
  output                                        mgr1__std__lane20_strm1_data_valid  ;

  input                                         std__mgr1__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane21_strm0_data        ;
  output                                        mgr1__std__lane21_strm0_data_valid  ;

  input                                         std__mgr1__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane21_strm1_data        ;
  output                                        mgr1__std__lane21_strm1_data_valid  ;

  input                                         std__mgr1__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane22_strm0_data        ;
  output                                        mgr1__std__lane22_strm0_data_valid  ;

  input                                         std__mgr1__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane22_strm1_data        ;
  output                                        mgr1__std__lane22_strm1_data_valid  ;

  input                                         std__mgr1__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane23_strm0_data        ;
  output                                        mgr1__std__lane23_strm0_data_valid  ;

  input                                         std__mgr1__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane23_strm1_data        ;
  output                                        mgr1__std__lane23_strm1_data_valid  ;

  input                                         std__mgr1__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane24_strm0_data        ;
  output                                        mgr1__std__lane24_strm0_data_valid  ;

  input                                         std__mgr1__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane24_strm1_data        ;
  output                                        mgr1__std__lane24_strm1_data_valid  ;

  input                                         std__mgr1__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane25_strm0_data        ;
  output                                        mgr1__std__lane25_strm0_data_valid  ;

  input                                         std__mgr1__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane25_strm1_data        ;
  output                                        mgr1__std__lane25_strm1_data_valid  ;

  input                                         std__mgr1__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane26_strm0_data        ;
  output                                        mgr1__std__lane26_strm0_data_valid  ;

  input                                         std__mgr1__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane26_strm1_data        ;
  output                                        mgr1__std__lane26_strm1_data_valid  ;

  input                                         std__mgr1__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane27_strm0_data        ;
  output                                        mgr1__std__lane27_strm0_data_valid  ;

  input                                         std__mgr1__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane27_strm1_data        ;
  output                                        mgr1__std__lane27_strm1_data_valid  ;

  input                                         std__mgr1__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane28_strm0_data        ;
  output                                        mgr1__std__lane28_strm0_data_valid  ;

  input                                         std__mgr1__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane28_strm1_data        ;
  output                                        mgr1__std__lane28_strm1_data_valid  ;

  input                                         std__mgr1__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane29_strm0_data        ;
  output                                        mgr1__std__lane29_strm0_data_valid  ;

  input                                         std__mgr1__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane29_strm1_data        ;
  output                                        mgr1__std__lane29_strm1_data_valid  ;

  input                                         std__mgr1__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane30_strm0_data        ;
  output                                        mgr1__std__lane30_strm0_data_valid  ;

  input                                         std__mgr1__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane30_strm1_data        ;
  output                                        mgr1__std__lane30_strm1_data_valid  ;

  input                                         std__mgr1__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane31_strm0_data        ;
  output                                        mgr1__std__lane31_strm0_data_valid  ;

  input                                         std__mgr1__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane31_strm1_data        ;
  output                                        mgr1__std__lane31_strm1_data_valid  ;

  input                                         std__mgr2__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane0_strm0_data        ;
  output                                        mgr2__std__lane0_strm0_data_valid  ;

  input                                         std__mgr2__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane0_strm1_data        ;
  output                                        mgr2__std__lane0_strm1_data_valid  ;

  input                                         std__mgr2__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane1_strm0_data        ;
  output                                        mgr2__std__lane1_strm0_data_valid  ;

  input                                         std__mgr2__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane1_strm1_data        ;
  output                                        mgr2__std__lane1_strm1_data_valid  ;

  input                                         std__mgr2__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane2_strm0_data        ;
  output                                        mgr2__std__lane2_strm0_data_valid  ;

  input                                         std__mgr2__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane2_strm1_data        ;
  output                                        mgr2__std__lane2_strm1_data_valid  ;

  input                                         std__mgr2__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane3_strm0_data        ;
  output                                        mgr2__std__lane3_strm0_data_valid  ;

  input                                         std__mgr2__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane3_strm1_data        ;
  output                                        mgr2__std__lane3_strm1_data_valid  ;

  input                                         std__mgr2__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane4_strm0_data        ;
  output                                        mgr2__std__lane4_strm0_data_valid  ;

  input                                         std__mgr2__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane4_strm1_data        ;
  output                                        mgr2__std__lane4_strm1_data_valid  ;

  input                                         std__mgr2__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane5_strm0_data        ;
  output                                        mgr2__std__lane5_strm0_data_valid  ;

  input                                         std__mgr2__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane5_strm1_data        ;
  output                                        mgr2__std__lane5_strm1_data_valid  ;

  input                                         std__mgr2__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane6_strm0_data        ;
  output                                        mgr2__std__lane6_strm0_data_valid  ;

  input                                         std__mgr2__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane6_strm1_data        ;
  output                                        mgr2__std__lane6_strm1_data_valid  ;

  input                                         std__mgr2__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane7_strm0_data        ;
  output                                        mgr2__std__lane7_strm0_data_valid  ;

  input                                         std__mgr2__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane7_strm1_data        ;
  output                                        mgr2__std__lane7_strm1_data_valid  ;

  input                                         std__mgr2__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane8_strm0_data        ;
  output                                        mgr2__std__lane8_strm0_data_valid  ;

  input                                         std__mgr2__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane8_strm1_data        ;
  output                                        mgr2__std__lane8_strm1_data_valid  ;

  input                                         std__mgr2__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane9_strm0_data        ;
  output                                        mgr2__std__lane9_strm0_data_valid  ;

  input                                         std__mgr2__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane9_strm1_data        ;
  output                                        mgr2__std__lane9_strm1_data_valid  ;

  input                                         std__mgr2__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane10_strm0_data        ;
  output                                        mgr2__std__lane10_strm0_data_valid  ;

  input                                         std__mgr2__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane10_strm1_data        ;
  output                                        mgr2__std__lane10_strm1_data_valid  ;

  input                                         std__mgr2__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane11_strm0_data        ;
  output                                        mgr2__std__lane11_strm0_data_valid  ;

  input                                         std__mgr2__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane11_strm1_data        ;
  output                                        mgr2__std__lane11_strm1_data_valid  ;

  input                                         std__mgr2__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane12_strm0_data        ;
  output                                        mgr2__std__lane12_strm0_data_valid  ;

  input                                         std__mgr2__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane12_strm1_data        ;
  output                                        mgr2__std__lane12_strm1_data_valid  ;

  input                                         std__mgr2__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane13_strm0_data        ;
  output                                        mgr2__std__lane13_strm0_data_valid  ;

  input                                         std__mgr2__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane13_strm1_data        ;
  output                                        mgr2__std__lane13_strm1_data_valid  ;

  input                                         std__mgr2__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane14_strm0_data        ;
  output                                        mgr2__std__lane14_strm0_data_valid  ;

  input                                         std__mgr2__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane14_strm1_data        ;
  output                                        mgr2__std__lane14_strm1_data_valid  ;

  input                                         std__mgr2__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane15_strm0_data        ;
  output                                        mgr2__std__lane15_strm0_data_valid  ;

  input                                         std__mgr2__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane15_strm1_data        ;
  output                                        mgr2__std__lane15_strm1_data_valid  ;

  input                                         std__mgr2__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane16_strm0_data        ;
  output                                        mgr2__std__lane16_strm0_data_valid  ;

  input                                         std__mgr2__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane16_strm1_data        ;
  output                                        mgr2__std__lane16_strm1_data_valid  ;

  input                                         std__mgr2__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane17_strm0_data        ;
  output                                        mgr2__std__lane17_strm0_data_valid  ;

  input                                         std__mgr2__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane17_strm1_data        ;
  output                                        mgr2__std__lane17_strm1_data_valid  ;

  input                                         std__mgr2__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane18_strm0_data        ;
  output                                        mgr2__std__lane18_strm0_data_valid  ;

  input                                         std__mgr2__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane18_strm1_data        ;
  output                                        mgr2__std__lane18_strm1_data_valid  ;

  input                                         std__mgr2__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane19_strm0_data        ;
  output                                        mgr2__std__lane19_strm0_data_valid  ;

  input                                         std__mgr2__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane19_strm1_data        ;
  output                                        mgr2__std__lane19_strm1_data_valid  ;

  input                                         std__mgr2__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane20_strm0_data        ;
  output                                        mgr2__std__lane20_strm0_data_valid  ;

  input                                         std__mgr2__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane20_strm1_data        ;
  output                                        mgr2__std__lane20_strm1_data_valid  ;

  input                                         std__mgr2__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane21_strm0_data        ;
  output                                        mgr2__std__lane21_strm0_data_valid  ;

  input                                         std__mgr2__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane21_strm1_data        ;
  output                                        mgr2__std__lane21_strm1_data_valid  ;

  input                                         std__mgr2__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane22_strm0_data        ;
  output                                        mgr2__std__lane22_strm0_data_valid  ;

  input                                         std__mgr2__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane22_strm1_data        ;
  output                                        mgr2__std__lane22_strm1_data_valid  ;

  input                                         std__mgr2__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane23_strm0_data        ;
  output                                        mgr2__std__lane23_strm0_data_valid  ;

  input                                         std__mgr2__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane23_strm1_data        ;
  output                                        mgr2__std__lane23_strm1_data_valid  ;

  input                                         std__mgr2__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane24_strm0_data        ;
  output                                        mgr2__std__lane24_strm0_data_valid  ;

  input                                         std__mgr2__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane24_strm1_data        ;
  output                                        mgr2__std__lane24_strm1_data_valid  ;

  input                                         std__mgr2__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane25_strm0_data        ;
  output                                        mgr2__std__lane25_strm0_data_valid  ;

  input                                         std__mgr2__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane25_strm1_data        ;
  output                                        mgr2__std__lane25_strm1_data_valid  ;

  input                                         std__mgr2__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane26_strm0_data        ;
  output                                        mgr2__std__lane26_strm0_data_valid  ;

  input                                         std__mgr2__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane26_strm1_data        ;
  output                                        mgr2__std__lane26_strm1_data_valid  ;

  input                                         std__mgr2__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane27_strm0_data        ;
  output                                        mgr2__std__lane27_strm0_data_valid  ;

  input                                         std__mgr2__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane27_strm1_data        ;
  output                                        mgr2__std__lane27_strm1_data_valid  ;

  input                                         std__mgr2__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane28_strm0_data        ;
  output                                        mgr2__std__lane28_strm0_data_valid  ;

  input                                         std__mgr2__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane28_strm1_data        ;
  output                                        mgr2__std__lane28_strm1_data_valid  ;

  input                                         std__mgr2__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane29_strm0_data        ;
  output                                        mgr2__std__lane29_strm0_data_valid  ;

  input                                         std__mgr2__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane29_strm1_data        ;
  output                                        mgr2__std__lane29_strm1_data_valid  ;

  input                                         std__mgr2__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane30_strm0_data        ;
  output                                        mgr2__std__lane30_strm0_data_valid  ;

  input                                         std__mgr2__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane30_strm1_data        ;
  output                                        mgr2__std__lane30_strm1_data_valid  ;

  input                                         std__mgr2__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane31_strm0_data        ;
  output                                        mgr2__std__lane31_strm0_data_valid  ;

  input                                         std__mgr2__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane31_strm1_data        ;
  output                                        mgr2__std__lane31_strm1_data_valid  ;

  input                                         std__mgr3__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane0_strm0_data        ;
  output                                        mgr3__std__lane0_strm0_data_valid  ;

  input                                         std__mgr3__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane0_strm1_data        ;
  output                                        mgr3__std__lane0_strm1_data_valid  ;

  input                                         std__mgr3__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane1_strm0_data        ;
  output                                        mgr3__std__lane1_strm0_data_valid  ;

  input                                         std__mgr3__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane1_strm1_data        ;
  output                                        mgr3__std__lane1_strm1_data_valid  ;

  input                                         std__mgr3__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane2_strm0_data        ;
  output                                        mgr3__std__lane2_strm0_data_valid  ;

  input                                         std__mgr3__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane2_strm1_data        ;
  output                                        mgr3__std__lane2_strm1_data_valid  ;

  input                                         std__mgr3__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane3_strm0_data        ;
  output                                        mgr3__std__lane3_strm0_data_valid  ;

  input                                         std__mgr3__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane3_strm1_data        ;
  output                                        mgr3__std__lane3_strm1_data_valid  ;

  input                                         std__mgr3__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane4_strm0_data        ;
  output                                        mgr3__std__lane4_strm0_data_valid  ;

  input                                         std__mgr3__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane4_strm1_data        ;
  output                                        mgr3__std__lane4_strm1_data_valid  ;

  input                                         std__mgr3__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane5_strm0_data        ;
  output                                        mgr3__std__lane5_strm0_data_valid  ;

  input                                         std__mgr3__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane5_strm1_data        ;
  output                                        mgr3__std__lane5_strm1_data_valid  ;

  input                                         std__mgr3__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane6_strm0_data        ;
  output                                        mgr3__std__lane6_strm0_data_valid  ;

  input                                         std__mgr3__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane6_strm1_data        ;
  output                                        mgr3__std__lane6_strm1_data_valid  ;

  input                                         std__mgr3__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane7_strm0_data        ;
  output                                        mgr3__std__lane7_strm0_data_valid  ;

  input                                         std__mgr3__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane7_strm1_data        ;
  output                                        mgr3__std__lane7_strm1_data_valid  ;

  input                                         std__mgr3__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane8_strm0_data        ;
  output                                        mgr3__std__lane8_strm0_data_valid  ;

  input                                         std__mgr3__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane8_strm1_data        ;
  output                                        mgr3__std__lane8_strm1_data_valid  ;

  input                                         std__mgr3__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane9_strm0_data        ;
  output                                        mgr3__std__lane9_strm0_data_valid  ;

  input                                         std__mgr3__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane9_strm1_data        ;
  output                                        mgr3__std__lane9_strm1_data_valid  ;

  input                                         std__mgr3__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane10_strm0_data        ;
  output                                        mgr3__std__lane10_strm0_data_valid  ;

  input                                         std__mgr3__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane10_strm1_data        ;
  output                                        mgr3__std__lane10_strm1_data_valid  ;

  input                                         std__mgr3__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane11_strm0_data        ;
  output                                        mgr3__std__lane11_strm0_data_valid  ;

  input                                         std__mgr3__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane11_strm1_data        ;
  output                                        mgr3__std__lane11_strm1_data_valid  ;

  input                                         std__mgr3__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane12_strm0_data        ;
  output                                        mgr3__std__lane12_strm0_data_valid  ;

  input                                         std__mgr3__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane12_strm1_data        ;
  output                                        mgr3__std__lane12_strm1_data_valid  ;

  input                                         std__mgr3__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane13_strm0_data        ;
  output                                        mgr3__std__lane13_strm0_data_valid  ;

  input                                         std__mgr3__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane13_strm1_data        ;
  output                                        mgr3__std__lane13_strm1_data_valid  ;

  input                                         std__mgr3__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane14_strm0_data        ;
  output                                        mgr3__std__lane14_strm0_data_valid  ;

  input                                         std__mgr3__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane14_strm1_data        ;
  output                                        mgr3__std__lane14_strm1_data_valid  ;

  input                                         std__mgr3__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane15_strm0_data        ;
  output                                        mgr3__std__lane15_strm0_data_valid  ;

  input                                         std__mgr3__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane15_strm1_data        ;
  output                                        mgr3__std__lane15_strm1_data_valid  ;

  input                                         std__mgr3__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane16_strm0_data        ;
  output                                        mgr3__std__lane16_strm0_data_valid  ;

  input                                         std__mgr3__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane16_strm1_data        ;
  output                                        mgr3__std__lane16_strm1_data_valid  ;

  input                                         std__mgr3__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane17_strm0_data        ;
  output                                        mgr3__std__lane17_strm0_data_valid  ;

  input                                         std__mgr3__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane17_strm1_data        ;
  output                                        mgr3__std__lane17_strm1_data_valid  ;

  input                                         std__mgr3__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane18_strm0_data        ;
  output                                        mgr3__std__lane18_strm0_data_valid  ;

  input                                         std__mgr3__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane18_strm1_data        ;
  output                                        mgr3__std__lane18_strm1_data_valid  ;

  input                                         std__mgr3__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane19_strm0_data        ;
  output                                        mgr3__std__lane19_strm0_data_valid  ;

  input                                         std__mgr3__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane19_strm1_data        ;
  output                                        mgr3__std__lane19_strm1_data_valid  ;

  input                                         std__mgr3__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane20_strm0_data        ;
  output                                        mgr3__std__lane20_strm0_data_valid  ;

  input                                         std__mgr3__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane20_strm1_data        ;
  output                                        mgr3__std__lane20_strm1_data_valid  ;

  input                                         std__mgr3__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane21_strm0_data        ;
  output                                        mgr3__std__lane21_strm0_data_valid  ;

  input                                         std__mgr3__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane21_strm1_data        ;
  output                                        mgr3__std__lane21_strm1_data_valid  ;

  input                                         std__mgr3__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane22_strm0_data        ;
  output                                        mgr3__std__lane22_strm0_data_valid  ;

  input                                         std__mgr3__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane22_strm1_data        ;
  output                                        mgr3__std__lane22_strm1_data_valid  ;

  input                                         std__mgr3__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane23_strm0_data        ;
  output                                        mgr3__std__lane23_strm0_data_valid  ;

  input                                         std__mgr3__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane23_strm1_data        ;
  output                                        mgr3__std__lane23_strm1_data_valid  ;

  input                                         std__mgr3__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane24_strm0_data        ;
  output                                        mgr3__std__lane24_strm0_data_valid  ;

  input                                         std__mgr3__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane24_strm1_data        ;
  output                                        mgr3__std__lane24_strm1_data_valid  ;

  input                                         std__mgr3__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane25_strm0_data        ;
  output                                        mgr3__std__lane25_strm0_data_valid  ;

  input                                         std__mgr3__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane25_strm1_data        ;
  output                                        mgr3__std__lane25_strm1_data_valid  ;

  input                                         std__mgr3__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane26_strm0_data        ;
  output                                        mgr3__std__lane26_strm0_data_valid  ;

  input                                         std__mgr3__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane26_strm1_data        ;
  output                                        mgr3__std__lane26_strm1_data_valid  ;

  input                                         std__mgr3__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane27_strm0_data        ;
  output                                        mgr3__std__lane27_strm0_data_valid  ;

  input                                         std__mgr3__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane27_strm1_data        ;
  output                                        mgr3__std__lane27_strm1_data_valid  ;

  input                                         std__mgr3__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane28_strm0_data        ;
  output                                        mgr3__std__lane28_strm0_data_valid  ;

  input                                         std__mgr3__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane28_strm1_data        ;
  output                                        mgr3__std__lane28_strm1_data_valid  ;

  input                                         std__mgr3__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane29_strm0_data        ;
  output                                        mgr3__std__lane29_strm0_data_valid  ;

  input                                         std__mgr3__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane29_strm1_data        ;
  output                                        mgr3__std__lane29_strm1_data_valid  ;

  input                                         std__mgr3__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane30_strm0_data        ;
  output                                        mgr3__std__lane30_strm0_data_valid  ;

  input                                         std__mgr3__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane30_strm1_data        ;
  output                                        mgr3__std__lane30_strm1_data_valid  ;

  input                                         std__mgr3__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane31_strm0_data        ;
  output                                        mgr3__std__lane31_strm0_data_valid  ;

  input                                         std__mgr3__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane31_strm1_data        ;
  output                                        mgr3__std__lane31_strm1_data_valid  ;

  input                                         std__mgr4__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane0_strm0_data        ;
  output                                        mgr4__std__lane0_strm0_data_valid  ;

  input                                         std__mgr4__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane0_strm1_data        ;
  output                                        mgr4__std__lane0_strm1_data_valid  ;

  input                                         std__mgr4__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane1_strm0_data        ;
  output                                        mgr4__std__lane1_strm0_data_valid  ;

  input                                         std__mgr4__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane1_strm1_data        ;
  output                                        mgr4__std__lane1_strm1_data_valid  ;

  input                                         std__mgr4__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane2_strm0_data        ;
  output                                        mgr4__std__lane2_strm0_data_valid  ;

  input                                         std__mgr4__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane2_strm1_data        ;
  output                                        mgr4__std__lane2_strm1_data_valid  ;

  input                                         std__mgr4__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane3_strm0_data        ;
  output                                        mgr4__std__lane3_strm0_data_valid  ;

  input                                         std__mgr4__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane3_strm1_data        ;
  output                                        mgr4__std__lane3_strm1_data_valid  ;

  input                                         std__mgr4__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane4_strm0_data        ;
  output                                        mgr4__std__lane4_strm0_data_valid  ;

  input                                         std__mgr4__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane4_strm1_data        ;
  output                                        mgr4__std__lane4_strm1_data_valid  ;

  input                                         std__mgr4__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane5_strm0_data        ;
  output                                        mgr4__std__lane5_strm0_data_valid  ;

  input                                         std__mgr4__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane5_strm1_data        ;
  output                                        mgr4__std__lane5_strm1_data_valid  ;

  input                                         std__mgr4__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane6_strm0_data        ;
  output                                        mgr4__std__lane6_strm0_data_valid  ;

  input                                         std__mgr4__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane6_strm1_data        ;
  output                                        mgr4__std__lane6_strm1_data_valid  ;

  input                                         std__mgr4__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane7_strm0_data        ;
  output                                        mgr4__std__lane7_strm0_data_valid  ;

  input                                         std__mgr4__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane7_strm1_data        ;
  output                                        mgr4__std__lane7_strm1_data_valid  ;

  input                                         std__mgr4__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane8_strm0_data        ;
  output                                        mgr4__std__lane8_strm0_data_valid  ;

  input                                         std__mgr4__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane8_strm1_data        ;
  output                                        mgr4__std__lane8_strm1_data_valid  ;

  input                                         std__mgr4__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane9_strm0_data        ;
  output                                        mgr4__std__lane9_strm0_data_valid  ;

  input                                         std__mgr4__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane9_strm1_data        ;
  output                                        mgr4__std__lane9_strm1_data_valid  ;

  input                                         std__mgr4__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane10_strm0_data        ;
  output                                        mgr4__std__lane10_strm0_data_valid  ;

  input                                         std__mgr4__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane10_strm1_data        ;
  output                                        mgr4__std__lane10_strm1_data_valid  ;

  input                                         std__mgr4__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane11_strm0_data        ;
  output                                        mgr4__std__lane11_strm0_data_valid  ;

  input                                         std__mgr4__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane11_strm1_data        ;
  output                                        mgr4__std__lane11_strm1_data_valid  ;

  input                                         std__mgr4__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane12_strm0_data        ;
  output                                        mgr4__std__lane12_strm0_data_valid  ;

  input                                         std__mgr4__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane12_strm1_data        ;
  output                                        mgr4__std__lane12_strm1_data_valid  ;

  input                                         std__mgr4__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane13_strm0_data        ;
  output                                        mgr4__std__lane13_strm0_data_valid  ;

  input                                         std__mgr4__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane13_strm1_data        ;
  output                                        mgr4__std__lane13_strm1_data_valid  ;

  input                                         std__mgr4__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane14_strm0_data        ;
  output                                        mgr4__std__lane14_strm0_data_valid  ;

  input                                         std__mgr4__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane14_strm1_data        ;
  output                                        mgr4__std__lane14_strm1_data_valid  ;

  input                                         std__mgr4__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane15_strm0_data        ;
  output                                        mgr4__std__lane15_strm0_data_valid  ;

  input                                         std__mgr4__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane15_strm1_data        ;
  output                                        mgr4__std__lane15_strm1_data_valid  ;

  input                                         std__mgr4__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane16_strm0_data        ;
  output                                        mgr4__std__lane16_strm0_data_valid  ;

  input                                         std__mgr4__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane16_strm1_data        ;
  output                                        mgr4__std__lane16_strm1_data_valid  ;

  input                                         std__mgr4__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane17_strm0_data        ;
  output                                        mgr4__std__lane17_strm0_data_valid  ;

  input                                         std__mgr4__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane17_strm1_data        ;
  output                                        mgr4__std__lane17_strm1_data_valid  ;

  input                                         std__mgr4__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane18_strm0_data        ;
  output                                        mgr4__std__lane18_strm0_data_valid  ;

  input                                         std__mgr4__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane18_strm1_data        ;
  output                                        mgr4__std__lane18_strm1_data_valid  ;

  input                                         std__mgr4__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane19_strm0_data        ;
  output                                        mgr4__std__lane19_strm0_data_valid  ;

  input                                         std__mgr4__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane19_strm1_data        ;
  output                                        mgr4__std__lane19_strm1_data_valid  ;

  input                                         std__mgr4__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane20_strm0_data        ;
  output                                        mgr4__std__lane20_strm0_data_valid  ;

  input                                         std__mgr4__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane20_strm1_data        ;
  output                                        mgr4__std__lane20_strm1_data_valid  ;

  input                                         std__mgr4__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane21_strm0_data        ;
  output                                        mgr4__std__lane21_strm0_data_valid  ;

  input                                         std__mgr4__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane21_strm1_data        ;
  output                                        mgr4__std__lane21_strm1_data_valid  ;

  input                                         std__mgr4__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane22_strm0_data        ;
  output                                        mgr4__std__lane22_strm0_data_valid  ;

  input                                         std__mgr4__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane22_strm1_data        ;
  output                                        mgr4__std__lane22_strm1_data_valid  ;

  input                                         std__mgr4__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane23_strm0_data        ;
  output                                        mgr4__std__lane23_strm0_data_valid  ;

  input                                         std__mgr4__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane23_strm1_data        ;
  output                                        mgr4__std__lane23_strm1_data_valid  ;

  input                                         std__mgr4__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane24_strm0_data        ;
  output                                        mgr4__std__lane24_strm0_data_valid  ;

  input                                         std__mgr4__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane24_strm1_data        ;
  output                                        mgr4__std__lane24_strm1_data_valid  ;

  input                                         std__mgr4__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane25_strm0_data        ;
  output                                        mgr4__std__lane25_strm0_data_valid  ;

  input                                         std__mgr4__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane25_strm1_data        ;
  output                                        mgr4__std__lane25_strm1_data_valid  ;

  input                                         std__mgr4__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane26_strm0_data        ;
  output                                        mgr4__std__lane26_strm0_data_valid  ;

  input                                         std__mgr4__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane26_strm1_data        ;
  output                                        mgr4__std__lane26_strm1_data_valid  ;

  input                                         std__mgr4__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane27_strm0_data        ;
  output                                        mgr4__std__lane27_strm0_data_valid  ;

  input                                         std__mgr4__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane27_strm1_data        ;
  output                                        mgr4__std__lane27_strm1_data_valid  ;

  input                                         std__mgr4__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane28_strm0_data        ;
  output                                        mgr4__std__lane28_strm0_data_valid  ;

  input                                         std__mgr4__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane28_strm1_data        ;
  output                                        mgr4__std__lane28_strm1_data_valid  ;

  input                                         std__mgr4__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane29_strm0_data        ;
  output                                        mgr4__std__lane29_strm0_data_valid  ;

  input                                         std__mgr4__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane29_strm1_data        ;
  output                                        mgr4__std__lane29_strm1_data_valid  ;

  input                                         std__mgr4__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane30_strm0_data        ;
  output                                        mgr4__std__lane30_strm0_data_valid  ;

  input                                         std__mgr4__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane30_strm1_data        ;
  output                                        mgr4__std__lane30_strm1_data_valid  ;

  input                                         std__mgr4__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane31_strm0_data        ;
  output                                        mgr4__std__lane31_strm0_data_valid  ;

  input                                         std__mgr4__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane31_strm1_data        ;
  output                                        mgr4__std__lane31_strm1_data_valid  ;

  input                                         std__mgr5__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane0_strm0_data        ;
  output                                        mgr5__std__lane0_strm0_data_valid  ;

  input                                         std__mgr5__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane0_strm1_data        ;
  output                                        mgr5__std__lane0_strm1_data_valid  ;

  input                                         std__mgr5__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane1_strm0_data        ;
  output                                        mgr5__std__lane1_strm0_data_valid  ;

  input                                         std__mgr5__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane1_strm1_data        ;
  output                                        mgr5__std__lane1_strm1_data_valid  ;

  input                                         std__mgr5__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane2_strm0_data        ;
  output                                        mgr5__std__lane2_strm0_data_valid  ;

  input                                         std__mgr5__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane2_strm1_data        ;
  output                                        mgr5__std__lane2_strm1_data_valid  ;

  input                                         std__mgr5__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane3_strm0_data        ;
  output                                        mgr5__std__lane3_strm0_data_valid  ;

  input                                         std__mgr5__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane3_strm1_data        ;
  output                                        mgr5__std__lane3_strm1_data_valid  ;

  input                                         std__mgr5__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane4_strm0_data        ;
  output                                        mgr5__std__lane4_strm0_data_valid  ;

  input                                         std__mgr5__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane4_strm1_data        ;
  output                                        mgr5__std__lane4_strm1_data_valid  ;

  input                                         std__mgr5__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane5_strm0_data        ;
  output                                        mgr5__std__lane5_strm0_data_valid  ;

  input                                         std__mgr5__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane5_strm1_data        ;
  output                                        mgr5__std__lane5_strm1_data_valid  ;

  input                                         std__mgr5__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane6_strm0_data        ;
  output                                        mgr5__std__lane6_strm0_data_valid  ;

  input                                         std__mgr5__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane6_strm1_data        ;
  output                                        mgr5__std__lane6_strm1_data_valid  ;

  input                                         std__mgr5__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane7_strm0_data        ;
  output                                        mgr5__std__lane7_strm0_data_valid  ;

  input                                         std__mgr5__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane7_strm1_data        ;
  output                                        mgr5__std__lane7_strm1_data_valid  ;

  input                                         std__mgr5__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane8_strm0_data        ;
  output                                        mgr5__std__lane8_strm0_data_valid  ;

  input                                         std__mgr5__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane8_strm1_data        ;
  output                                        mgr5__std__lane8_strm1_data_valid  ;

  input                                         std__mgr5__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane9_strm0_data        ;
  output                                        mgr5__std__lane9_strm0_data_valid  ;

  input                                         std__mgr5__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane9_strm1_data        ;
  output                                        mgr5__std__lane9_strm1_data_valid  ;

  input                                         std__mgr5__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane10_strm0_data        ;
  output                                        mgr5__std__lane10_strm0_data_valid  ;

  input                                         std__mgr5__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane10_strm1_data        ;
  output                                        mgr5__std__lane10_strm1_data_valid  ;

  input                                         std__mgr5__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane11_strm0_data        ;
  output                                        mgr5__std__lane11_strm0_data_valid  ;

  input                                         std__mgr5__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane11_strm1_data        ;
  output                                        mgr5__std__lane11_strm1_data_valid  ;

  input                                         std__mgr5__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane12_strm0_data        ;
  output                                        mgr5__std__lane12_strm0_data_valid  ;

  input                                         std__mgr5__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane12_strm1_data        ;
  output                                        mgr5__std__lane12_strm1_data_valid  ;

  input                                         std__mgr5__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane13_strm0_data        ;
  output                                        mgr5__std__lane13_strm0_data_valid  ;

  input                                         std__mgr5__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane13_strm1_data        ;
  output                                        mgr5__std__lane13_strm1_data_valid  ;

  input                                         std__mgr5__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane14_strm0_data        ;
  output                                        mgr5__std__lane14_strm0_data_valid  ;

  input                                         std__mgr5__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane14_strm1_data        ;
  output                                        mgr5__std__lane14_strm1_data_valid  ;

  input                                         std__mgr5__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane15_strm0_data        ;
  output                                        mgr5__std__lane15_strm0_data_valid  ;

  input                                         std__mgr5__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane15_strm1_data        ;
  output                                        mgr5__std__lane15_strm1_data_valid  ;

  input                                         std__mgr5__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane16_strm0_data        ;
  output                                        mgr5__std__lane16_strm0_data_valid  ;

  input                                         std__mgr5__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane16_strm1_data        ;
  output                                        mgr5__std__lane16_strm1_data_valid  ;

  input                                         std__mgr5__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane17_strm0_data        ;
  output                                        mgr5__std__lane17_strm0_data_valid  ;

  input                                         std__mgr5__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane17_strm1_data        ;
  output                                        mgr5__std__lane17_strm1_data_valid  ;

  input                                         std__mgr5__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane18_strm0_data        ;
  output                                        mgr5__std__lane18_strm0_data_valid  ;

  input                                         std__mgr5__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane18_strm1_data        ;
  output                                        mgr5__std__lane18_strm1_data_valid  ;

  input                                         std__mgr5__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane19_strm0_data        ;
  output                                        mgr5__std__lane19_strm0_data_valid  ;

  input                                         std__mgr5__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane19_strm1_data        ;
  output                                        mgr5__std__lane19_strm1_data_valid  ;

  input                                         std__mgr5__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane20_strm0_data        ;
  output                                        mgr5__std__lane20_strm0_data_valid  ;

  input                                         std__mgr5__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane20_strm1_data        ;
  output                                        mgr5__std__lane20_strm1_data_valid  ;

  input                                         std__mgr5__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane21_strm0_data        ;
  output                                        mgr5__std__lane21_strm0_data_valid  ;

  input                                         std__mgr5__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane21_strm1_data        ;
  output                                        mgr5__std__lane21_strm1_data_valid  ;

  input                                         std__mgr5__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane22_strm0_data        ;
  output                                        mgr5__std__lane22_strm0_data_valid  ;

  input                                         std__mgr5__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane22_strm1_data        ;
  output                                        mgr5__std__lane22_strm1_data_valid  ;

  input                                         std__mgr5__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane23_strm0_data        ;
  output                                        mgr5__std__lane23_strm0_data_valid  ;

  input                                         std__mgr5__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane23_strm1_data        ;
  output                                        mgr5__std__lane23_strm1_data_valid  ;

  input                                         std__mgr5__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane24_strm0_data        ;
  output                                        mgr5__std__lane24_strm0_data_valid  ;

  input                                         std__mgr5__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane24_strm1_data        ;
  output                                        mgr5__std__lane24_strm1_data_valid  ;

  input                                         std__mgr5__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane25_strm0_data        ;
  output                                        mgr5__std__lane25_strm0_data_valid  ;

  input                                         std__mgr5__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane25_strm1_data        ;
  output                                        mgr5__std__lane25_strm1_data_valid  ;

  input                                         std__mgr5__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane26_strm0_data        ;
  output                                        mgr5__std__lane26_strm0_data_valid  ;

  input                                         std__mgr5__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane26_strm1_data        ;
  output                                        mgr5__std__lane26_strm1_data_valid  ;

  input                                         std__mgr5__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane27_strm0_data        ;
  output                                        mgr5__std__lane27_strm0_data_valid  ;

  input                                         std__mgr5__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane27_strm1_data        ;
  output                                        mgr5__std__lane27_strm1_data_valid  ;

  input                                         std__mgr5__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane28_strm0_data        ;
  output                                        mgr5__std__lane28_strm0_data_valid  ;

  input                                         std__mgr5__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane28_strm1_data        ;
  output                                        mgr5__std__lane28_strm1_data_valid  ;

  input                                         std__mgr5__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane29_strm0_data        ;
  output                                        mgr5__std__lane29_strm0_data_valid  ;

  input                                         std__mgr5__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane29_strm1_data        ;
  output                                        mgr5__std__lane29_strm1_data_valid  ;

  input                                         std__mgr5__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane30_strm0_data        ;
  output                                        mgr5__std__lane30_strm0_data_valid  ;

  input                                         std__mgr5__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane30_strm1_data        ;
  output                                        mgr5__std__lane30_strm1_data_valid  ;

  input                                         std__mgr5__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane31_strm0_data        ;
  output                                        mgr5__std__lane31_strm0_data_valid  ;

  input                                         std__mgr5__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane31_strm1_data        ;
  output                                        mgr5__std__lane31_strm1_data_valid  ;

  input                                         std__mgr6__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane0_strm0_data        ;
  output                                        mgr6__std__lane0_strm0_data_valid  ;

  input                                         std__mgr6__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane0_strm1_data        ;
  output                                        mgr6__std__lane0_strm1_data_valid  ;

  input                                         std__mgr6__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane1_strm0_data        ;
  output                                        mgr6__std__lane1_strm0_data_valid  ;

  input                                         std__mgr6__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane1_strm1_data        ;
  output                                        mgr6__std__lane1_strm1_data_valid  ;

  input                                         std__mgr6__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane2_strm0_data        ;
  output                                        mgr6__std__lane2_strm0_data_valid  ;

  input                                         std__mgr6__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane2_strm1_data        ;
  output                                        mgr6__std__lane2_strm1_data_valid  ;

  input                                         std__mgr6__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane3_strm0_data        ;
  output                                        mgr6__std__lane3_strm0_data_valid  ;

  input                                         std__mgr6__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane3_strm1_data        ;
  output                                        mgr6__std__lane3_strm1_data_valid  ;

  input                                         std__mgr6__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane4_strm0_data        ;
  output                                        mgr6__std__lane4_strm0_data_valid  ;

  input                                         std__mgr6__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane4_strm1_data        ;
  output                                        mgr6__std__lane4_strm1_data_valid  ;

  input                                         std__mgr6__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane5_strm0_data        ;
  output                                        mgr6__std__lane5_strm0_data_valid  ;

  input                                         std__mgr6__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane5_strm1_data        ;
  output                                        mgr6__std__lane5_strm1_data_valid  ;

  input                                         std__mgr6__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane6_strm0_data        ;
  output                                        mgr6__std__lane6_strm0_data_valid  ;

  input                                         std__mgr6__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane6_strm1_data        ;
  output                                        mgr6__std__lane6_strm1_data_valid  ;

  input                                         std__mgr6__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane7_strm0_data        ;
  output                                        mgr6__std__lane7_strm0_data_valid  ;

  input                                         std__mgr6__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane7_strm1_data        ;
  output                                        mgr6__std__lane7_strm1_data_valid  ;

  input                                         std__mgr6__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane8_strm0_data        ;
  output                                        mgr6__std__lane8_strm0_data_valid  ;

  input                                         std__mgr6__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane8_strm1_data        ;
  output                                        mgr6__std__lane8_strm1_data_valid  ;

  input                                         std__mgr6__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane9_strm0_data        ;
  output                                        mgr6__std__lane9_strm0_data_valid  ;

  input                                         std__mgr6__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane9_strm1_data        ;
  output                                        mgr6__std__lane9_strm1_data_valid  ;

  input                                         std__mgr6__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane10_strm0_data        ;
  output                                        mgr6__std__lane10_strm0_data_valid  ;

  input                                         std__mgr6__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane10_strm1_data        ;
  output                                        mgr6__std__lane10_strm1_data_valid  ;

  input                                         std__mgr6__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane11_strm0_data        ;
  output                                        mgr6__std__lane11_strm0_data_valid  ;

  input                                         std__mgr6__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane11_strm1_data        ;
  output                                        mgr6__std__lane11_strm1_data_valid  ;

  input                                         std__mgr6__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane12_strm0_data        ;
  output                                        mgr6__std__lane12_strm0_data_valid  ;

  input                                         std__mgr6__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane12_strm1_data        ;
  output                                        mgr6__std__lane12_strm1_data_valid  ;

  input                                         std__mgr6__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane13_strm0_data        ;
  output                                        mgr6__std__lane13_strm0_data_valid  ;

  input                                         std__mgr6__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane13_strm1_data        ;
  output                                        mgr6__std__lane13_strm1_data_valid  ;

  input                                         std__mgr6__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane14_strm0_data        ;
  output                                        mgr6__std__lane14_strm0_data_valid  ;

  input                                         std__mgr6__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane14_strm1_data        ;
  output                                        mgr6__std__lane14_strm1_data_valid  ;

  input                                         std__mgr6__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane15_strm0_data        ;
  output                                        mgr6__std__lane15_strm0_data_valid  ;

  input                                         std__mgr6__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane15_strm1_data        ;
  output                                        mgr6__std__lane15_strm1_data_valid  ;

  input                                         std__mgr6__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane16_strm0_data        ;
  output                                        mgr6__std__lane16_strm0_data_valid  ;

  input                                         std__mgr6__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane16_strm1_data        ;
  output                                        mgr6__std__lane16_strm1_data_valid  ;

  input                                         std__mgr6__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane17_strm0_data        ;
  output                                        mgr6__std__lane17_strm0_data_valid  ;

  input                                         std__mgr6__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane17_strm1_data        ;
  output                                        mgr6__std__lane17_strm1_data_valid  ;

  input                                         std__mgr6__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane18_strm0_data        ;
  output                                        mgr6__std__lane18_strm0_data_valid  ;

  input                                         std__mgr6__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane18_strm1_data        ;
  output                                        mgr6__std__lane18_strm1_data_valid  ;

  input                                         std__mgr6__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane19_strm0_data        ;
  output                                        mgr6__std__lane19_strm0_data_valid  ;

  input                                         std__mgr6__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane19_strm1_data        ;
  output                                        mgr6__std__lane19_strm1_data_valid  ;

  input                                         std__mgr6__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane20_strm0_data        ;
  output                                        mgr6__std__lane20_strm0_data_valid  ;

  input                                         std__mgr6__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane20_strm1_data        ;
  output                                        mgr6__std__lane20_strm1_data_valid  ;

  input                                         std__mgr6__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane21_strm0_data        ;
  output                                        mgr6__std__lane21_strm0_data_valid  ;

  input                                         std__mgr6__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane21_strm1_data        ;
  output                                        mgr6__std__lane21_strm1_data_valid  ;

  input                                         std__mgr6__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane22_strm0_data        ;
  output                                        mgr6__std__lane22_strm0_data_valid  ;

  input                                         std__mgr6__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane22_strm1_data        ;
  output                                        mgr6__std__lane22_strm1_data_valid  ;

  input                                         std__mgr6__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane23_strm0_data        ;
  output                                        mgr6__std__lane23_strm0_data_valid  ;

  input                                         std__mgr6__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane23_strm1_data        ;
  output                                        mgr6__std__lane23_strm1_data_valid  ;

  input                                         std__mgr6__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane24_strm0_data        ;
  output                                        mgr6__std__lane24_strm0_data_valid  ;

  input                                         std__mgr6__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane24_strm1_data        ;
  output                                        mgr6__std__lane24_strm1_data_valid  ;

  input                                         std__mgr6__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane25_strm0_data        ;
  output                                        mgr6__std__lane25_strm0_data_valid  ;

  input                                         std__mgr6__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane25_strm1_data        ;
  output                                        mgr6__std__lane25_strm1_data_valid  ;

  input                                         std__mgr6__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane26_strm0_data        ;
  output                                        mgr6__std__lane26_strm0_data_valid  ;

  input                                         std__mgr6__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane26_strm1_data        ;
  output                                        mgr6__std__lane26_strm1_data_valid  ;

  input                                         std__mgr6__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane27_strm0_data        ;
  output                                        mgr6__std__lane27_strm0_data_valid  ;

  input                                         std__mgr6__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane27_strm1_data        ;
  output                                        mgr6__std__lane27_strm1_data_valid  ;

  input                                         std__mgr6__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane28_strm0_data        ;
  output                                        mgr6__std__lane28_strm0_data_valid  ;

  input                                         std__mgr6__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane28_strm1_data        ;
  output                                        mgr6__std__lane28_strm1_data_valid  ;

  input                                         std__mgr6__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane29_strm0_data        ;
  output                                        mgr6__std__lane29_strm0_data_valid  ;

  input                                         std__mgr6__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane29_strm1_data        ;
  output                                        mgr6__std__lane29_strm1_data_valid  ;

  input                                         std__mgr6__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane30_strm0_data        ;
  output                                        mgr6__std__lane30_strm0_data_valid  ;

  input                                         std__mgr6__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane30_strm1_data        ;
  output                                        mgr6__std__lane30_strm1_data_valid  ;

  input                                         std__mgr6__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane31_strm0_data        ;
  output                                        mgr6__std__lane31_strm0_data_valid  ;

  input                                         std__mgr6__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane31_strm1_data        ;
  output                                        mgr6__std__lane31_strm1_data_valid  ;

  input                                         std__mgr7__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane0_strm0_data        ;
  output                                        mgr7__std__lane0_strm0_data_valid  ;

  input                                         std__mgr7__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane0_strm1_data        ;
  output                                        mgr7__std__lane0_strm1_data_valid  ;

  input                                         std__mgr7__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane1_strm0_data        ;
  output                                        mgr7__std__lane1_strm0_data_valid  ;

  input                                         std__mgr7__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane1_strm1_data        ;
  output                                        mgr7__std__lane1_strm1_data_valid  ;

  input                                         std__mgr7__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane2_strm0_data        ;
  output                                        mgr7__std__lane2_strm0_data_valid  ;

  input                                         std__mgr7__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane2_strm1_data        ;
  output                                        mgr7__std__lane2_strm1_data_valid  ;

  input                                         std__mgr7__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane3_strm0_data        ;
  output                                        mgr7__std__lane3_strm0_data_valid  ;

  input                                         std__mgr7__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane3_strm1_data        ;
  output                                        mgr7__std__lane3_strm1_data_valid  ;

  input                                         std__mgr7__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane4_strm0_data        ;
  output                                        mgr7__std__lane4_strm0_data_valid  ;

  input                                         std__mgr7__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane4_strm1_data        ;
  output                                        mgr7__std__lane4_strm1_data_valid  ;

  input                                         std__mgr7__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane5_strm0_data        ;
  output                                        mgr7__std__lane5_strm0_data_valid  ;

  input                                         std__mgr7__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane5_strm1_data        ;
  output                                        mgr7__std__lane5_strm1_data_valid  ;

  input                                         std__mgr7__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane6_strm0_data        ;
  output                                        mgr7__std__lane6_strm0_data_valid  ;

  input                                         std__mgr7__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane6_strm1_data        ;
  output                                        mgr7__std__lane6_strm1_data_valid  ;

  input                                         std__mgr7__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane7_strm0_data        ;
  output                                        mgr7__std__lane7_strm0_data_valid  ;

  input                                         std__mgr7__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane7_strm1_data        ;
  output                                        mgr7__std__lane7_strm1_data_valid  ;

  input                                         std__mgr7__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane8_strm0_data        ;
  output                                        mgr7__std__lane8_strm0_data_valid  ;

  input                                         std__mgr7__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane8_strm1_data        ;
  output                                        mgr7__std__lane8_strm1_data_valid  ;

  input                                         std__mgr7__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane9_strm0_data        ;
  output                                        mgr7__std__lane9_strm0_data_valid  ;

  input                                         std__mgr7__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane9_strm1_data        ;
  output                                        mgr7__std__lane9_strm1_data_valid  ;

  input                                         std__mgr7__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane10_strm0_data        ;
  output                                        mgr7__std__lane10_strm0_data_valid  ;

  input                                         std__mgr7__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane10_strm1_data        ;
  output                                        mgr7__std__lane10_strm1_data_valid  ;

  input                                         std__mgr7__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane11_strm0_data        ;
  output                                        mgr7__std__lane11_strm0_data_valid  ;

  input                                         std__mgr7__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane11_strm1_data        ;
  output                                        mgr7__std__lane11_strm1_data_valid  ;

  input                                         std__mgr7__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane12_strm0_data        ;
  output                                        mgr7__std__lane12_strm0_data_valid  ;

  input                                         std__mgr7__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane12_strm1_data        ;
  output                                        mgr7__std__lane12_strm1_data_valid  ;

  input                                         std__mgr7__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane13_strm0_data        ;
  output                                        mgr7__std__lane13_strm0_data_valid  ;

  input                                         std__mgr7__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane13_strm1_data        ;
  output                                        mgr7__std__lane13_strm1_data_valid  ;

  input                                         std__mgr7__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane14_strm0_data        ;
  output                                        mgr7__std__lane14_strm0_data_valid  ;

  input                                         std__mgr7__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane14_strm1_data        ;
  output                                        mgr7__std__lane14_strm1_data_valid  ;

  input                                         std__mgr7__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane15_strm0_data        ;
  output                                        mgr7__std__lane15_strm0_data_valid  ;

  input                                         std__mgr7__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane15_strm1_data        ;
  output                                        mgr7__std__lane15_strm1_data_valid  ;

  input                                         std__mgr7__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane16_strm0_data        ;
  output                                        mgr7__std__lane16_strm0_data_valid  ;

  input                                         std__mgr7__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane16_strm1_data        ;
  output                                        mgr7__std__lane16_strm1_data_valid  ;

  input                                         std__mgr7__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane17_strm0_data        ;
  output                                        mgr7__std__lane17_strm0_data_valid  ;

  input                                         std__mgr7__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane17_strm1_data        ;
  output                                        mgr7__std__lane17_strm1_data_valid  ;

  input                                         std__mgr7__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane18_strm0_data        ;
  output                                        mgr7__std__lane18_strm0_data_valid  ;

  input                                         std__mgr7__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane18_strm1_data        ;
  output                                        mgr7__std__lane18_strm1_data_valid  ;

  input                                         std__mgr7__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane19_strm0_data        ;
  output                                        mgr7__std__lane19_strm0_data_valid  ;

  input                                         std__mgr7__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane19_strm1_data        ;
  output                                        mgr7__std__lane19_strm1_data_valid  ;

  input                                         std__mgr7__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane20_strm0_data        ;
  output                                        mgr7__std__lane20_strm0_data_valid  ;

  input                                         std__mgr7__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane20_strm1_data        ;
  output                                        mgr7__std__lane20_strm1_data_valid  ;

  input                                         std__mgr7__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane21_strm0_data        ;
  output                                        mgr7__std__lane21_strm0_data_valid  ;

  input                                         std__mgr7__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane21_strm1_data        ;
  output                                        mgr7__std__lane21_strm1_data_valid  ;

  input                                         std__mgr7__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane22_strm0_data        ;
  output                                        mgr7__std__lane22_strm0_data_valid  ;

  input                                         std__mgr7__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane22_strm1_data        ;
  output                                        mgr7__std__lane22_strm1_data_valid  ;

  input                                         std__mgr7__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane23_strm0_data        ;
  output                                        mgr7__std__lane23_strm0_data_valid  ;

  input                                         std__mgr7__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane23_strm1_data        ;
  output                                        mgr7__std__lane23_strm1_data_valid  ;

  input                                         std__mgr7__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane24_strm0_data        ;
  output                                        mgr7__std__lane24_strm0_data_valid  ;

  input                                         std__mgr7__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane24_strm1_data        ;
  output                                        mgr7__std__lane24_strm1_data_valid  ;

  input                                         std__mgr7__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane25_strm0_data        ;
  output                                        mgr7__std__lane25_strm0_data_valid  ;

  input                                         std__mgr7__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane25_strm1_data        ;
  output                                        mgr7__std__lane25_strm1_data_valid  ;

  input                                         std__mgr7__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane26_strm0_data        ;
  output                                        mgr7__std__lane26_strm0_data_valid  ;

  input                                         std__mgr7__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane26_strm1_data        ;
  output                                        mgr7__std__lane26_strm1_data_valid  ;

  input                                         std__mgr7__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane27_strm0_data        ;
  output                                        mgr7__std__lane27_strm0_data_valid  ;

  input                                         std__mgr7__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane27_strm1_data        ;
  output                                        mgr7__std__lane27_strm1_data_valid  ;

  input                                         std__mgr7__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane28_strm0_data        ;
  output                                        mgr7__std__lane28_strm0_data_valid  ;

  input                                         std__mgr7__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane28_strm1_data        ;
  output                                        mgr7__std__lane28_strm1_data_valid  ;

  input                                         std__mgr7__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane29_strm0_data        ;
  output                                        mgr7__std__lane29_strm0_data_valid  ;

  input                                         std__mgr7__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane29_strm1_data        ;
  output                                        mgr7__std__lane29_strm1_data_valid  ;

  input                                         std__mgr7__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane30_strm0_data        ;
  output                                        mgr7__std__lane30_strm0_data_valid  ;

  input                                         std__mgr7__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane30_strm1_data        ;
  output                                        mgr7__std__lane30_strm1_data_valid  ;

  input                                         std__mgr7__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane31_strm0_data        ;
  output                                        mgr7__std__lane31_strm0_data_valid  ;

  input                                         std__mgr7__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane31_strm1_data        ;
  output                                        mgr7__std__lane31_strm1_data_valid  ;

  input                                         std__mgr8__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane0_strm0_data        ;
  output                                        mgr8__std__lane0_strm0_data_valid  ;

  input                                         std__mgr8__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane0_strm1_data        ;
  output                                        mgr8__std__lane0_strm1_data_valid  ;

  input                                         std__mgr8__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane1_strm0_data        ;
  output                                        mgr8__std__lane1_strm0_data_valid  ;

  input                                         std__mgr8__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane1_strm1_data        ;
  output                                        mgr8__std__lane1_strm1_data_valid  ;

  input                                         std__mgr8__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane2_strm0_data        ;
  output                                        mgr8__std__lane2_strm0_data_valid  ;

  input                                         std__mgr8__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane2_strm1_data        ;
  output                                        mgr8__std__lane2_strm1_data_valid  ;

  input                                         std__mgr8__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane3_strm0_data        ;
  output                                        mgr8__std__lane3_strm0_data_valid  ;

  input                                         std__mgr8__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane3_strm1_data        ;
  output                                        mgr8__std__lane3_strm1_data_valid  ;

  input                                         std__mgr8__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane4_strm0_data        ;
  output                                        mgr8__std__lane4_strm0_data_valid  ;

  input                                         std__mgr8__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane4_strm1_data        ;
  output                                        mgr8__std__lane4_strm1_data_valid  ;

  input                                         std__mgr8__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane5_strm0_data        ;
  output                                        mgr8__std__lane5_strm0_data_valid  ;

  input                                         std__mgr8__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane5_strm1_data        ;
  output                                        mgr8__std__lane5_strm1_data_valid  ;

  input                                         std__mgr8__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane6_strm0_data        ;
  output                                        mgr8__std__lane6_strm0_data_valid  ;

  input                                         std__mgr8__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane6_strm1_data        ;
  output                                        mgr8__std__lane6_strm1_data_valid  ;

  input                                         std__mgr8__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane7_strm0_data        ;
  output                                        mgr8__std__lane7_strm0_data_valid  ;

  input                                         std__mgr8__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane7_strm1_data        ;
  output                                        mgr8__std__lane7_strm1_data_valid  ;

  input                                         std__mgr8__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane8_strm0_data        ;
  output                                        mgr8__std__lane8_strm0_data_valid  ;

  input                                         std__mgr8__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane8_strm1_data        ;
  output                                        mgr8__std__lane8_strm1_data_valid  ;

  input                                         std__mgr8__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane9_strm0_data        ;
  output                                        mgr8__std__lane9_strm0_data_valid  ;

  input                                         std__mgr8__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane9_strm1_data        ;
  output                                        mgr8__std__lane9_strm1_data_valid  ;

  input                                         std__mgr8__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane10_strm0_data        ;
  output                                        mgr8__std__lane10_strm0_data_valid  ;

  input                                         std__mgr8__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane10_strm1_data        ;
  output                                        mgr8__std__lane10_strm1_data_valid  ;

  input                                         std__mgr8__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane11_strm0_data        ;
  output                                        mgr8__std__lane11_strm0_data_valid  ;

  input                                         std__mgr8__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane11_strm1_data        ;
  output                                        mgr8__std__lane11_strm1_data_valid  ;

  input                                         std__mgr8__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane12_strm0_data        ;
  output                                        mgr8__std__lane12_strm0_data_valid  ;

  input                                         std__mgr8__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane12_strm1_data        ;
  output                                        mgr8__std__lane12_strm1_data_valid  ;

  input                                         std__mgr8__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane13_strm0_data        ;
  output                                        mgr8__std__lane13_strm0_data_valid  ;

  input                                         std__mgr8__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane13_strm1_data        ;
  output                                        mgr8__std__lane13_strm1_data_valid  ;

  input                                         std__mgr8__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane14_strm0_data        ;
  output                                        mgr8__std__lane14_strm0_data_valid  ;

  input                                         std__mgr8__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane14_strm1_data        ;
  output                                        mgr8__std__lane14_strm1_data_valid  ;

  input                                         std__mgr8__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane15_strm0_data        ;
  output                                        mgr8__std__lane15_strm0_data_valid  ;

  input                                         std__mgr8__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane15_strm1_data        ;
  output                                        mgr8__std__lane15_strm1_data_valid  ;

  input                                         std__mgr8__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane16_strm0_data        ;
  output                                        mgr8__std__lane16_strm0_data_valid  ;

  input                                         std__mgr8__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane16_strm1_data        ;
  output                                        mgr8__std__lane16_strm1_data_valid  ;

  input                                         std__mgr8__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane17_strm0_data        ;
  output                                        mgr8__std__lane17_strm0_data_valid  ;

  input                                         std__mgr8__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane17_strm1_data        ;
  output                                        mgr8__std__lane17_strm1_data_valid  ;

  input                                         std__mgr8__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane18_strm0_data        ;
  output                                        mgr8__std__lane18_strm0_data_valid  ;

  input                                         std__mgr8__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane18_strm1_data        ;
  output                                        mgr8__std__lane18_strm1_data_valid  ;

  input                                         std__mgr8__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane19_strm0_data        ;
  output                                        mgr8__std__lane19_strm0_data_valid  ;

  input                                         std__mgr8__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane19_strm1_data        ;
  output                                        mgr8__std__lane19_strm1_data_valid  ;

  input                                         std__mgr8__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane20_strm0_data        ;
  output                                        mgr8__std__lane20_strm0_data_valid  ;

  input                                         std__mgr8__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane20_strm1_data        ;
  output                                        mgr8__std__lane20_strm1_data_valid  ;

  input                                         std__mgr8__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane21_strm0_data        ;
  output                                        mgr8__std__lane21_strm0_data_valid  ;

  input                                         std__mgr8__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane21_strm1_data        ;
  output                                        mgr8__std__lane21_strm1_data_valid  ;

  input                                         std__mgr8__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane22_strm0_data        ;
  output                                        mgr8__std__lane22_strm0_data_valid  ;

  input                                         std__mgr8__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane22_strm1_data        ;
  output                                        mgr8__std__lane22_strm1_data_valid  ;

  input                                         std__mgr8__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane23_strm0_data        ;
  output                                        mgr8__std__lane23_strm0_data_valid  ;

  input                                         std__mgr8__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane23_strm1_data        ;
  output                                        mgr8__std__lane23_strm1_data_valid  ;

  input                                         std__mgr8__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane24_strm0_data        ;
  output                                        mgr8__std__lane24_strm0_data_valid  ;

  input                                         std__mgr8__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane24_strm1_data        ;
  output                                        mgr8__std__lane24_strm1_data_valid  ;

  input                                         std__mgr8__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane25_strm0_data        ;
  output                                        mgr8__std__lane25_strm0_data_valid  ;

  input                                         std__mgr8__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane25_strm1_data        ;
  output                                        mgr8__std__lane25_strm1_data_valid  ;

  input                                         std__mgr8__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane26_strm0_data        ;
  output                                        mgr8__std__lane26_strm0_data_valid  ;

  input                                         std__mgr8__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane26_strm1_data        ;
  output                                        mgr8__std__lane26_strm1_data_valid  ;

  input                                         std__mgr8__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane27_strm0_data        ;
  output                                        mgr8__std__lane27_strm0_data_valid  ;

  input                                         std__mgr8__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane27_strm1_data        ;
  output                                        mgr8__std__lane27_strm1_data_valid  ;

  input                                         std__mgr8__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane28_strm0_data        ;
  output                                        mgr8__std__lane28_strm0_data_valid  ;

  input                                         std__mgr8__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane28_strm1_data        ;
  output                                        mgr8__std__lane28_strm1_data_valid  ;

  input                                         std__mgr8__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane29_strm0_data        ;
  output                                        mgr8__std__lane29_strm0_data_valid  ;

  input                                         std__mgr8__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane29_strm1_data        ;
  output                                        mgr8__std__lane29_strm1_data_valid  ;

  input                                         std__mgr8__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane30_strm0_data        ;
  output                                        mgr8__std__lane30_strm0_data_valid  ;

  input                                         std__mgr8__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane30_strm1_data        ;
  output                                        mgr8__std__lane30_strm1_data_valid  ;

  input                                         std__mgr8__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane31_strm0_data        ;
  output                                        mgr8__std__lane31_strm0_data_valid  ;

  input                                         std__mgr8__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane31_strm1_data        ;
  output                                        mgr8__std__lane31_strm1_data_valid  ;

  input                                         std__mgr9__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane0_strm0_data        ;
  output                                        mgr9__std__lane0_strm0_data_valid  ;

  input                                         std__mgr9__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane0_strm1_data        ;
  output                                        mgr9__std__lane0_strm1_data_valid  ;

  input                                         std__mgr9__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane1_strm0_data        ;
  output                                        mgr9__std__lane1_strm0_data_valid  ;

  input                                         std__mgr9__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane1_strm1_data        ;
  output                                        mgr9__std__lane1_strm1_data_valid  ;

  input                                         std__mgr9__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane2_strm0_data        ;
  output                                        mgr9__std__lane2_strm0_data_valid  ;

  input                                         std__mgr9__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane2_strm1_data        ;
  output                                        mgr9__std__lane2_strm1_data_valid  ;

  input                                         std__mgr9__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane3_strm0_data        ;
  output                                        mgr9__std__lane3_strm0_data_valid  ;

  input                                         std__mgr9__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane3_strm1_data        ;
  output                                        mgr9__std__lane3_strm1_data_valid  ;

  input                                         std__mgr9__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane4_strm0_data        ;
  output                                        mgr9__std__lane4_strm0_data_valid  ;

  input                                         std__mgr9__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane4_strm1_data        ;
  output                                        mgr9__std__lane4_strm1_data_valid  ;

  input                                         std__mgr9__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane5_strm0_data        ;
  output                                        mgr9__std__lane5_strm0_data_valid  ;

  input                                         std__mgr9__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane5_strm1_data        ;
  output                                        mgr9__std__lane5_strm1_data_valid  ;

  input                                         std__mgr9__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane6_strm0_data        ;
  output                                        mgr9__std__lane6_strm0_data_valid  ;

  input                                         std__mgr9__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane6_strm1_data        ;
  output                                        mgr9__std__lane6_strm1_data_valid  ;

  input                                         std__mgr9__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane7_strm0_data        ;
  output                                        mgr9__std__lane7_strm0_data_valid  ;

  input                                         std__mgr9__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane7_strm1_data        ;
  output                                        mgr9__std__lane7_strm1_data_valid  ;

  input                                         std__mgr9__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane8_strm0_data        ;
  output                                        mgr9__std__lane8_strm0_data_valid  ;

  input                                         std__mgr9__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane8_strm1_data        ;
  output                                        mgr9__std__lane8_strm1_data_valid  ;

  input                                         std__mgr9__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane9_strm0_data        ;
  output                                        mgr9__std__lane9_strm0_data_valid  ;

  input                                         std__mgr9__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane9_strm1_data        ;
  output                                        mgr9__std__lane9_strm1_data_valid  ;

  input                                         std__mgr9__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane10_strm0_data        ;
  output                                        mgr9__std__lane10_strm0_data_valid  ;

  input                                         std__mgr9__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane10_strm1_data        ;
  output                                        mgr9__std__lane10_strm1_data_valid  ;

  input                                         std__mgr9__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane11_strm0_data        ;
  output                                        mgr9__std__lane11_strm0_data_valid  ;

  input                                         std__mgr9__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane11_strm1_data        ;
  output                                        mgr9__std__lane11_strm1_data_valid  ;

  input                                         std__mgr9__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane12_strm0_data        ;
  output                                        mgr9__std__lane12_strm0_data_valid  ;

  input                                         std__mgr9__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane12_strm1_data        ;
  output                                        mgr9__std__lane12_strm1_data_valid  ;

  input                                         std__mgr9__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane13_strm0_data        ;
  output                                        mgr9__std__lane13_strm0_data_valid  ;

  input                                         std__mgr9__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane13_strm1_data        ;
  output                                        mgr9__std__lane13_strm1_data_valid  ;

  input                                         std__mgr9__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane14_strm0_data        ;
  output                                        mgr9__std__lane14_strm0_data_valid  ;

  input                                         std__mgr9__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane14_strm1_data        ;
  output                                        mgr9__std__lane14_strm1_data_valid  ;

  input                                         std__mgr9__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane15_strm0_data        ;
  output                                        mgr9__std__lane15_strm0_data_valid  ;

  input                                         std__mgr9__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane15_strm1_data        ;
  output                                        mgr9__std__lane15_strm1_data_valid  ;

  input                                         std__mgr9__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane16_strm0_data        ;
  output                                        mgr9__std__lane16_strm0_data_valid  ;

  input                                         std__mgr9__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane16_strm1_data        ;
  output                                        mgr9__std__lane16_strm1_data_valid  ;

  input                                         std__mgr9__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane17_strm0_data        ;
  output                                        mgr9__std__lane17_strm0_data_valid  ;

  input                                         std__mgr9__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane17_strm1_data        ;
  output                                        mgr9__std__lane17_strm1_data_valid  ;

  input                                         std__mgr9__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane18_strm0_data        ;
  output                                        mgr9__std__lane18_strm0_data_valid  ;

  input                                         std__mgr9__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane18_strm1_data        ;
  output                                        mgr9__std__lane18_strm1_data_valid  ;

  input                                         std__mgr9__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane19_strm0_data        ;
  output                                        mgr9__std__lane19_strm0_data_valid  ;

  input                                         std__mgr9__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane19_strm1_data        ;
  output                                        mgr9__std__lane19_strm1_data_valid  ;

  input                                         std__mgr9__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane20_strm0_data        ;
  output                                        mgr9__std__lane20_strm0_data_valid  ;

  input                                         std__mgr9__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane20_strm1_data        ;
  output                                        mgr9__std__lane20_strm1_data_valid  ;

  input                                         std__mgr9__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane21_strm0_data        ;
  output                                        mgr9__std__lane21_strm0_data_valid  ;

  input                                         std__mgr9__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane21_strm1_data        ;
  output                                        mgr9__std__lane21_strm1_data_valid  ;

  input                                         std__mgr9__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane22_strm0_data        ;
  output                                        mgr9__std__lane22_strm0_data_valid  ;

  input                                         std__mgr9__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane22_strm1_data        ;
  output                                        mgr9__std__lane22_strm1_data_valid  ;

  input                                         std__mgr9__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane23_strm0_data        ;
  output                                        mgr9__std__lane23_strm0_data_valid  ;

  input                                         std__mgr9__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane23_strm1_data        ;
  output                                        mgr9__std__lane23_strm1_data_valid  ;

  input                                         std__mgr9__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane24_strm0_data        ;
  output                                        mgr9__std__lane24_strm0_data_valid  ;

  input                                         std__mgr9__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane24_strm1_data        ;
  output                                        mgr9__std__lane24_strm1_data_valid  ;

  input                                         std__mgr9__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane25_strm0_data        ;
  output                                        mgr9__std__lane25_strm0_data_valid  ;

  input                                         std__mgr9__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane25_strm1_data        ;
  output                                        mgr9__std__lane25_strm1_data_valid  ;

  input                                         std__mgr9__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane26_strm0_data        ;
  output                                        mgr9__std__lane26_strm0_data_valid  ;

  input                                         std__mgr9__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane26_strm1_data        ;
  output                                        mgr9__std__lane26_strm1_data_valid  ;

  input                                         std__mgr9__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane27_strm0_data        ;
  output                                        mgr9__std__lane27_strm0_data_valid  ;

  input                                         std__mgr9__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane27_strm1_data        ;
  output                                        mgr9__std__lane27_strm1_data_valid  ;

  input                                         std__mgr9__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane28_strm0_data        ;
  output                                        mgr9__std__lane28_strm0_data_valid  ;

  input                                         std__mgr9__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane28_strm1_data        ;
  output                                        mgr9__std__lane28_strm1_data_valid  ;

  input                                         std__mgr9__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane29_strm0_data        ;
  output                                        mgr9__std__lane29_strm0_data_valid  ;

  input                                         std__mgr9__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane29_strm1_data        ;
  output                                        mgr9__std__lane29_strm1_data_valid  ;

  input                                         std__mgr9__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane30_strm0_data        ;
  output                                        mgr9__std__lane30_strm0_data_valid  ;

  input                                         std__mgr9__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane30_strm1_data        ;
  output                                        mgr9__std__lane30_strm1_data_valid  ;

  input                                         std__mgr9__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane31_strm0_data        ;
  output                                        mgr9__std__lane31_strm0_data_valid  ;

  input                                         std__mgr9__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane31_strm1_data        ;
  output                                        mgr9__std__lane31_strm1_data_valid  ;

  input                                         std__mgr10__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane0_strm0_data        ;
  output                                        mgr10__std__lane0_strm0_data_valid  ;

  input                                         std__mgr10__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane0_strm1_data        ;
  output                                        mgr10__std__lane0_strm1_data_valid  ;

  input                                         std__mgr10__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane1_strm0_data        ;
  output                                        mgr10__std__lane1_strm0_data_valid  ;

  input                                         std__mgr10__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane1_strm1_data        ;
  output                                        mgr10__std__lane1_strm1_data_valid  ;

  input                                         std__mgr10__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane2_strm0_data        ;
  output                                        mgr10__std__lane2_strm0_data_valid  ;

  input                                         std__mgr10__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane2_strm1_data        ;
  output                                        mgr10__std__lane2_strm1_data_valid  ;

  input                                         std__mgr10__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane3_strm0_data        ;
  output                                        mgr10__std__lane3_strm0_data_valid  ;

  input                                         std__mgr10__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane3_strm1_data        ;
  output                                        mgr10__std__lane3_strm1_data_valid  ;

  input                                         std__mgr10__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane4_strm0_data        ;
  output                                        mgr10__std__lane4_strm0_data_valid  ;

  input                                         std__mgr10__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane4_strm1_data        ;
  output                                        mgr10__std__lane4_strm1_data_valid  ;

  input                                         std__mgr10__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane5_strm0_data        ;
  output                                        mgr10__std__lane5_strm0_data_valid  ;

  input                                         std__mgr10__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane5_strm1_data        ;
  output                                        mgr10__std__lane5_strm1_data_valid  ;

  input                                         std__mgr10__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane6_strm0_data        ;
  output                                        mgr10__std__lane6_strm0_data_valid  ;

  input                                         std__mgr10__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane6_strm1_data        ;
  output                                        mgr10__std__lane6_strm1_data_valid  ;

  input                                         std__mgr10__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane7_strm0_data        ;
  output                                        mgr10__std__lane7_strm0_data_valid  ;

  input                                         std__mgr10__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane7_strm1_data        ;
  output                                        mgr10__std__lane7_strm1_data_valid  ;

  input                                         std__mgr10__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane8_strm0_data        ;
  output                                        mgr10__std__lane8_strm0_data_valid  ;

  input                                         std__mgr10__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane8_strm1_data        ;
  output                                        mgr10__std__lane8_strm1_data_valid  ;

  input                                         std__mgr10__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane9_strm0_data        ;
  output                                        mgr10__std__lane9_strm0_data_valid  ;

  input                                         std__mgr10__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane9_strm1_data        ;
  output                                        mgr10__std__lane9_strm1_data_valid  ;

  input                                         std__mgr10__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane10_strm0_data        ;
  output                                        mgr10__std__lane10_strm0_data_valid  ;

  input                                         std__mgr10__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane10_strm1_data        ;
  output                                        mgr10__std__lane10_strm1_data_valid  ;

  input                                         std__mgr10__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane11_strm0_data        ;
  output                                        mgr10__std__lane11_strm0_data_valid  ;

  input                                         std__mgr10__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane11_strm1_data        ;
  output                                        mgr10__std__lane11_strm1_data_valid  ;

  input                                         std__mgr10__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane12_strm0_data        ;
  output                                        mgr10__std__lane12_strm0_data_valid  ;

  input                                         std__mgr10__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane12_strm1_data        ;
  output                                        mgr10__std__lane12_strm1_data_valid  ;

  input                                         std__mgr10__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane13_strm0_data        ;
  output                                        mgr10__std__lane13_strm0_data_valid  ;

  input                                         std__mgr10__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane13_strm1_data        ;
  output                                        mgr10__std__lane13_strm1_data_valid  ;

  input                                         std__mgr10__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane14_strm0_data        ;
  output                                        mgr10__std__lane14_strm0_data_valid  ;

  input                                         std__mgr10__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane14_strm1_data        ;
  output                                        mgr10__std__lane14_strm1_data_valid  ;

  input                                         std__mgr10__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane15_strm0_data        ;
  output                                        mgr10__std__lane15_strm0_data_valid  ;

  input                                         std__mgr10__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane15_strm1_data        ;
  output                                        mgr10__std__lane15_strm1_data_valid  ;

  input                                         std__mgr10__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane16_strm0_data        ;
  output                                        mgr10__std__lane16_strm0_data_valid  ;

  input                                         std__mgr10__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane16_strm1_data        ;
  output                                        mgr10__std__lane16_strm1_data_valid  ;

  input                                         std__mgr10__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane17_strm0_data        ;
  output                                        mgr10__std__lane17_strm0_data_valid  ;

  input                                         std__mgr10__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane17_strm1_data        ;
  output                                        mgr10__std__lane17_strm1_data_valid  ;

  input                                         std__mgr10__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane18_strm0_data        ;
  output                                        mgr10__std__lane18_strm0_data_valid  ;

  input                                         std__mgr10__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane18_strm1_data        ;
  output                                        mgr10__std__lane18_strm1_data_valid  ;

  input                                         std__mgr10__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane19_strm0_data        ;
  output                                        mgr10__std__lane19_strm0_data_valid  ;

  input                                         std__mgr10__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane19_strm1_data        ;
  output                                        mgr10__std__lane19_strm1_data_valid  ;

  input                                         std__mgr10__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane20_strm0_data        ;
  output                                        mgr10__std__lane20_strm0_data_valid  ;

  input                                         std__mgr10__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane20_strm1_data        ;
  output                                        mgr10__std__lane20_strm1_data_valid  ;

  input                                         std__mgr10__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane21_strm0_data        ;
  output                                        mgr10__std__lane21_strm0_data_valid  ;

  input                                         std__mgr10__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane21_strm1_data        ;
  output                                        mgr10__std__lane21_strm1_data_valid  ;

  input                                         std__mgr10__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane22_strm0_data        ;
  output                                        mgr10__std__lane22_strm0_data_valid  ;

  input                                         std__mgr10__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane22_strm1_data        ;
  output                                        mgr10__std__lane22_strm1_data_valid  ;

  input                                         std__mgr10__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane23_strm0_data        ;
  output                                        mgr10__std__lane23_strm0_data_valid  ;

  input                                         std__mgr10__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane23_strm1_data        ;
  output                                        mgr10__std__lane23_strm1_data_valid  ;

  input                                         std__mgr10__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane24_strm0_data        ;
  output                                        mgr10__std__lane24_strm0_data_valid  ;

  input                                         std__mgr10__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane24_strm1_data        ;
  output                                        mgr10__std__lane24_strm1_data_valid  ;

  input                                         std__mgr10__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane25_strm0_data        ;
  output                                        mgr10__std__lane25_strm0_data_valid  ;

  input                                         std__mgr10__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane25_strm1_data        ;
  output                                        mgr10__std__lane25_strm1_data_valid  ;

  input                                         std__mgr10__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane26_strm0_data        ;
  output                                        mgr10__std__lane26_strm0_data_valid  ;

  input                                         std__mgr10__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane26_strm1_data        ;
  output                                        mgr10__std__lane26_strm1_data_valid  ;

  input                                         std__mgr10__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane27_strm0_data        ;
  output                                        mgr10__std__lane27_strm0_data_valid  ;

  input                                         std__mgr10__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane27_strm1_data        ;
  output                                        mgr10__std__lane27_strm1_data_valid  ;

  input                                         std__mgr10__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane28_strm0_data        ;
  output                                        mgr10__std__lane28_strm0_data_valid  ;

  input                                         std__mgr10__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane28_strm1_data        ;
  output                                        mgr10__std__lane28_strm1_data_valid  ;

  input                                         std__mgr10__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane29_strm0_data        ;
  output                                        mgr10__std__lane29_strm0_data_valid  ;

  input                                         std__mgr10__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane29_strm1_data        ;
  output                                        mgr10__std__lane29_strm1_data_valid  ;

  input                                         std__mgr10__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane30_strm0_data        ;
  output                                        mgr10__std__lane30_strm0_data_valid  ;

  input                                         std__mgr10__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane30_strm1_data        ;
  output                                        mgr10__std__lane30_strm1_data_valid  ;

  input                                         std__mgr10__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane31_strm0_data        ;
  output                                        mgr10__std__lane31_strm0_data_valid  ;

  input                                         std__mgr10__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane31_strm1_data        ;
  output                                        mgr10__std__lane31_strm1_data_valid  ;

  input                                         std__mgr11__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane0_strm0_data        ;
  output                                        mgr11__std__lane0_strm0_data_valid  ;

  input                                         std__mgr11__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane0_strm1_data        ;
  output                                        mgr11__std__lane0_strm1_data_valid  ;

  input                                         std__mgr11__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane1_strm0_data        ;
  output                                        mgr11__std__lane1_strm0_data_valid  ;

  input                                         std__mgr11__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane1_strm1_data        ;
  output                                        mgr11__std__lane1_strm1_data_valid  ;

  input                                         std__mgr11__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane2_strm0_data        ;
  output                                        mgr11__std__lane2_strm0_data_valid  ;

  input                                         std__mgr11__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane2_strm1_data        ;
  output                                        mgr11__std__lane2_strm1_data_valid  ;

  input                                         std__mgr11__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane3_strm0_data        ;
  output                                        mgr11__std__lane3_strm0_data_valid  ;

  input                                         std__mgr11__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane3_strm1_data        ;
  output                                        mgr11__std__lane3_strm1_data_valid  ;

  input                                         std__mgr11__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane4_strm0_data        ;
  output                                        mgr11__std__lane4_strm0_data_valid  ;

  input                                         std__mgr11__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane4_strm1_data        ;
  output                                        mgr11__std__lane4_strm1_data_valid  ;

  input                                         std__mgr11__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane5_strm0_data        ;
  output                                        mgr11__std__lane5_strm0_data_valid  ;

  input                                         std__mgr11__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane5_strm1_data        ;
  output                                        mgr11__std__lane5_strm1_data_valid  ;

  input                                         std__mgr11__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane6_strm0_data        ;
  output                                        mgr11__std__lane6_strm0_data_valid  ;

  input                                         std__mgr11__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane6_strm1_data        ;
  output                                        mgr11__std__lane6_strm1_data_valid  ;

  input                                         std__mgr11__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane7_strm0_data        ;
  output                                        mgr11__std__lane7_strm0_data_valid  ;

  input                                         std__mgr11__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane7_strm1_data        ;
  output                                        mgr11__std__lane7_strm1_data_valid  ;

  input                                         std__mgr11__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane8_strm0_data        ;
  output                                        mgr11__std__lane8_strm0_data_valid  ;

  input                                         std__mgr11__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane8_strm1_data        ;
  output                                        mgr11__std__lane8_strm1_data_valid  ;

  input                                         std__mgr11__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane9_strm0_data        ;
  output                                        mgr11__std__lane9_strm0_data_valid  ;

  input                                         std__mgr11__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane9_strm1_data        ;
  output                                        mgr11__std__lane9_strm1_data_valid  ;

  input                                         std__mgr11__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane10_strm0_data        ;
  output                                        mgr11__std__lane10_strm0_data_valid  ;

  input                                         std__mgr11__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane10_strm1_data        ;
  output                                        mgr11__std__lane10_strm1_data_valid  ;

  input                                         std__mgr11__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane11_strm0_data        ;
  output                                        mgr11__std__lane11_strm0_data_valid  ;

  input                                         std__mgr11__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane11_strm1_data        ;
  output                                        mgr11__std__lane11_strm1_data_valid  ;

  input                                         std__mgr11__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane12_strm0_data        ;
  output                                        mgr11__std__lane12_strm0_data_valid  ;

  input                                         std__mgr11__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane12_strm1_data        ;
  output                                        mgr11__std__lane12_strm1_data_valid  ;

  input                                         std__mgr11__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane13_strm0_data        ;
  output                                        mgr11__std__lane13_strm0_data_valid  ;

  input                                         std__mgr11__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane13_strm1_data        ;
  output                                        mgr11__std__lane13_strm1_data_valid  ;

  input                                         std__mgr11__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane14_strm0_data        ;
  output                                        mgr11__std__lane14_strm0_data_valid  ;

  input                                         std__mgr11__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane14_strm1_data        ;
  output                                        mgr11__std__lane14_strm1_data_valid  ;

  input                                         std__mgr11__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane15_strm0_data        ;
  output                                        mgr11__std__lane15_strm0_data_valid  ;

  input                                         std__mgr11__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane15_strm1_data        ;
  output                                        mgr11__std__lane15_strm1_data_valid  ;

  input                                         std__mgr11__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane16_strm0_data        ;
  output                                        mgr11__std__lane16_strm0_data_valid  ;

  input                                         std__mgr11__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane16_strm1_data        ;
  output                                        mgr11__std__lane16_strm1_data_valid  ;

  input                                         std__mgr11__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane17_strm0_data        ;
  output                                        mgr11__std__lane17_strm0_data_valid  ;

  input                                         std__mgr11__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane17_strm1_data        ;
  output                                        mgr11__std__lane17_strm1_data_valid  ;

  input                                         std__mgr11__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane18_strm0_data        ;
  output                                        mgr11__std__lane18_strm0_data_valid  ;

  input                                         std__mgr11__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane18_strm1_data        ;
  output                                        mgr11__std__lane18_strm1_data_valid  ;

  input                                         std__mgr11__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane19_strm0_data        ;
  output                                        mgr11__std__lane19_strm0_data_valid  ;

  input                                         std__mgr11__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane19_strm1_data        ;
  output                                        mgr11__std__lane19_strm1_data_valid  ;

  input                                         std__mgr11__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane20_strm0_data        ;
  output                                        mgr11__std__lane20_strm0_data_valid  ;

  input                                         std__mgr11__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane20_strm1_data        ;
  output                                        mgr11__std__lane20_strm1_data_valid  ;

  input                                         std__mgr11__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane21_strm0_data        ;
  output                                        mgr11__std__lane21_strm0_data_valid  ;

  input                                         std__mgr11__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane21_strm1_data        ;
  output                                        mgr11__std__lane21_strm1_data_valid  ;

  input                                         std__mgr11__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane22_strm0_data        ;
  output                                        mgr11__std__lane22_strm0_data_valid  ;

  input                                         std__mgr11__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane22_strm1_data        ;
  output                                        mgr11__std__lane22_strm1_data_valid  ;

  input                                         std__mgr11__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane23_strm0_data        ;
  output                                        mgr11__std__lane23_strm0_data_valid  ;

  input                                         std__mgr11__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane23_strm1_data        ;
  output                                        mgr11__std__lane23_strm1_data_valid  ;

  input                                         std__mgr11__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane24_strm0_data        ;
  output                                        mgr11__std__lane24_strm0_data_valid  ;

  input                                         std__mgr11__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane24_strm1_data        ;
  output                                        mgr11__std__lane24_strm1_data_valid  ;

  input                                         std__mgr11__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane25_strm0_data        ;
  output                                        mgr11__std__lane25_strm0_data_valid  ;

  input                                         std__mgr11__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane25_strm1_data        ;
  output                                        mgr11__std__lane25_strm1_data_valid  ;

  input                                         std__mgr11__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane26_strm0_data        ;
  output                                        mgr11__std__lane26_strm0_data_valid  ;

  input                                         std__mgr11__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane26_strm1_data        ;
  output                                        mgr11__std__lane26_strm1_data_valid  ;

  input                                         std__mgr11__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane27_strm0_data        ;
  output                                        mgr11__std__lane27_strm0_data_valid  ;

  input                                         std__mgr11__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane27_strm1_data        ;
  output                                        mgr11__std__lane27_strm1_data_valid  ;

  input                                         std__mgr11__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane28_strm0_data        ;
  output                                        mgr11__std__lane28_strm0_data_valid  ;

  input                                         std__mgr11__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane28_strm1_data        ;
  output                                        mgr11__std__lane28_strm1_data_valid  ;

  input                                         std__mgr11__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane29_strm0_data        ;
  output                                        mgr11__std__lane29_strm0_data_valid  ;

  input                                         std__mgr11__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane29_strm1_data        ;
  output                                        mgr11__std__lane29_strm1_data_valid  ;

  input                                         std__mgr11__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane30_strm0_data        ;
  output                                        mgr11__std__lane30_strm0_data_valid  ;

  input                                         std__mgr11__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane30_strm1_data        ;
  output                                        mgr11__std__lane30_strm1_data_valid  ;

  input                                         std__mgr11__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane31_strm0_data        ;
  output                                        mgr11__std__lane31_strm0_data_valid  ;

  input                                         std__mgr11__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane31_strm1_data        ;
  output                                        mgr11__std__lane31_strm1_data_valid  ;

  input                                         std__mgr12__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane0_strm0_data        ;
  output                                        mgr12__std__lane0_strm0_data_valid  ;

  input                                         std__mgr12__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane0_strm1_data        ;
  output                                        mgr12__std__lane0_strm1_data_valid  ;

  input                                         std__mgr12__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane1_strm0_data        ;
  output                                        mgr12__std__lane1_strm0_data_valid  ;

  input                                         std__mgr12__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane1_strm1_data        ;
  output                                        mgr12__std__lane1_strm1_data_valid  ;

  input                                         std__mgr12__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane2_strm0_data        ;
  output                                        mgr12__std__lane2_strm0_data_valid  ;

  input                                         std__mgr12__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane2_strm1_data        ;
  output                                        mgr12__std__lane2_strm1_data_valid  ;

  input                                         std__mgr12__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane3_strm0_data        ;
  output                                        mgr12__std__lane3_strm0_data_valid  ;

  input                                         std__mgr12__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane3_strm1_data        ;
  output                                        mgr12__std__lane3_strm1_data_valid  ;

  input                                         std__mgr12__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane4_strm0_data        ;
  output                                        mgr12__std__lane4_strm0_data_valid  ;

  input                                         std__mgr12__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane4_strm1_data        ;
  output                                        mgr12__std__lane4_strm1_data_valid  ;

  input                                         std__mgr12__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane5_strm0_data        ;
  output                                        mgr12__std__lane5_strm0_data_valid  ;

  input                                         std__mgr12__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane5_strm1_data        ;
  output                                        mgr12__std__lane5_strm1_data_valid  ;

  input                                         std__mgr12__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane6_strm0_data        ;
  output                                        mgr12__std__lane6_strm0_data_valid  ;

  input                                         std__mgr12__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane6_strm1_data        ;
  output                                        mgr12__std__lane6_strm1_data_valid  ;

  input                                         std__mgr12__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane7_strm0_data        ;
  output                                        mgr12__std__lane7_strm0_data_valid  ;

  input                                         std__mgr12__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane7_strm1_data        ;
  output                                        mgr12__std__lane7_strm1_data_valid  ;

  input                                         std__mgr12__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane8_strm0_data        ;
  output                                        mgr12__std__lane8_strm0_data_valid  ;

  input                                         std__mgr12__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane8_strm1_data        ;
  output                                        mgr12__std__lane8_strm1_data_valid  ;

  input                                         std__mgr12__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane9_strm0_data        ;
  output                                        mgr12__std__lane9_strm0_data_valid  ;

  input                                         std__mgr12__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane9_strm1_data        ;
  output                                        mgr12__std__lane9_strm1_data_valid  ;

  input                                         std__mgr12__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane10_strm0_data        ;
  output                                        mgr12__std__lane10_strm0_data_valid  ;

  input                                         std__mgr12__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane10_strm1_data        ;
  output                                        mgr12__std__lane10_strm1_data_valid  ;

  input                                         std__mgr12__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane11_strm0_data        ;
  output                                        mgr12__std__lane11_strm0_data_valid  ;

  input                                         std__mgr12__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane11_strm1_data        ;
  output                                        mgr12__std__lane11_strm1_data_valid  ;

  input                                         std__mgr12__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane12_strm0_data        ;
  output                                        mgr12__std__lane12_strm0_data_valid  ;

  input                                         std__mgr12__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane12_strm1_data        ;
  output                                        mgr12__std__lane12_strm1_data_valid  ;

  input                                         std__mgr12__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane13_strm0_data        ;
  output                                        mgr12__std__lane13_strm0_data_valid  ;

  input                                         std__mgr12__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane13_strm1_data        ;
  output                                        mgr12__std__lane13_strm1_data_valid  ;

  input                                         std__mgr12__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane14_strm0_data        ;
  output                                        mgr12__std__lane14_strm0_data_valid  ;

  input                                         std__mgr12__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane14_strm1_data        ;
  output                                        mgr12__std__lane14_strm1_data_valid  ;

  input                                         std__mgr12__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane15_strm0_data        ;
  output                                        mgr12__std__lane15_strm0_data_valid  ;

  input                                         std__mgr12__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane15_strm1_data        ;
  output                                        mgr12__std__lane15_strm1_data_valid  ;

  input                                         std__mgr12__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane16_strm0_data        ;
  output                                        mgr12__std__lane16_strm0_data_valid  ;

  input                                         std__mgr12__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane16_strm1_data        ;
  output                                        mgr12__std__lane16_strm1_data_valid  ;

  input                                         std__mgr12__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane17_strm0_data        ;
  output                                        mgr12__std__lane17_strm0_data_valid  ;

  input                                         std__mgr12__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane17_strm1_data        ;
  output                                        mgr12__std__lane17_strm1_data_valid  ;

  input                                         std__mgr12__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane18_strm0_data        ;
  output                                        mgr12__std__lane18_strm0_data_valid  ;

  input                                         std__mgr12__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane18_strm1_data        ;
  output                                        mgr12__std__lane18_strm1_data_valid  ;

  input                                         std__mgr12__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane19_strm0_data        ;
  output                                        mgr12__std__lane19_strm0_data_valid  ;

  input                                         std__mgr12__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane19_strm1_data        ;
  output                                        mgr12__std__lane19_strm1_data_valid  ;

  input                                         std__mgr12__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane20_strm0_data        ;
  output                                        mgr12__std__lane20_strm0_data_valid  ;

  input                                         std__mgr12__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane20_strm1_data        ;
  output                                        mgr12__std__lane20_strm1_data_valid  ;

  input                                         std__mgr12__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane21_strm0_data        ;
  output                                        mgr12__std__lane21_strm0_data_valid  ;

  input                                         std__mgr12__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane21_strm1_data        ;
  output                                        mgr12__std__lane21_strm1_data_valid  ;

  input                                         std__mgr12__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane22_strm0_data        ;
  output                                        mgr12__std__lane22_strm0_data_valid  ;

  input                                         std__mgr12__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane22_strm1_data        ;
  output                                        mgr12__std__lane22_strm1_data_valid  ;

  input                                         std__mgr12__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane23_strm0_data        ;
  output                                        mgr12__std__lane23_strm0_data_valid  ;

  input                                         std__mgr12__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane23_strm1_data        ;
  output                                        mgr12__std__lane23_strm1_data_valid  ;

  input                                         std__mgr12__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane24_strm0_data        ;
  output                                        mgr12__std__lane24_strm0_data_valid  ;

  input                                         std__mgr12__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane24_strm1_data        ;
  output                                        mgr12__std__lane24_strm1_data_valid  ;

  input                                         std__mgr12__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane25_strm0_data        ;
  output                                        mgr12__std__lane25_strm0_data_valid  ;

  input                                         std__mgr12__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane25_strm1_data        ;
  output                                        mgr12__std__lane25_strm1_data_valid  ;

  input                                         std__mgr12__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane26_strm0_data        ;
  output                                        mgr12__std__lane26_strm0_data_valid  ;

  input                                         std__mgr12__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane26_strm1_data        ;
  output                                        mgr12__std__lane26_strm1_data_valid  ;

  input                                         std__mgr12__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane27_strm0_data        ;
  output                                        mgr12__std__lane27_strm0_data_valid  ;

  input                                         std__mgr12__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane27_strm1_data        ;
  output                                        mgr12__std__lane27_strm1_data_valid  ;

  input                                         std__mgr12__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane28_strm0_data        ;
  output                                        mgr12__std__lane28_strm0_data_valid  ;

  input                                         std__mgr12__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane28_strm1_data        ;
  output                                        mgr12__std__lane28_strm1_data_valid  ;

  input                                         std__mgr12__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane29_strm0_data        ;
  output                                        mgr12__std__lane29_strm0_data_valid  ;

  input                                         std__mgr12__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane29_strm1_data        ;
  output                                        mgr12__std__lane29_strm1_data_valid  ;

  input                                         std__mgr12__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane30_strm0_data        ;
  output                                        mgr12__std__lane30_strm0_data_valid  ;

  input                                         std__mgr12__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane30_strm1_data        ;
  output                                        mgr12__std__lane30_strm1_data_valid  ;

  input                                         std__mgr12__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane31_strm0_data        ;
  output                                        mgr12__std__lane31_strm0_data_valid  ;

  input                                         std__mgr12__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane31_strm1_data        ;
  output                                        mgr12__std__lane31_strm1_data_valid  ;

  input                                         std__mgr13__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane0_strm0_data        ;
  output                                        mgr13__std__lane0_strm0_data_valid  ;

  input                                         std__mgr13__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane0_strm1_data        ;
  output                                        mgr13__std__lane0_strm1_data_valid  ;

  input                                         std__mgr13__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane1_strm0_data        ;
  output                                        mgr13__std__lane1_strm0_data_valid  ;

  input                                         std__mgr13__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane1_strm1_data        ;
  output                                        mgr13__std__lane1_strm1_data_valid  ;

  input                                         std__mgr13__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane2_strm0_data        ;
  output                                        mgr13__std__lane2_strm0_data_valid  ;

  input                                         std__mgr13__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane2_strm1_data        ;
  output                                        mgr13__std__lane2_strm1_data_valid  ;

  input                                         std__mgr13__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane3_strm0_data        ;
  output                                        mgr13__std__lane3_strm0_data_valid  ;

  input                                         std__mgr13__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane3_strm1_data        ;
  output                                        mgr13__std__lane3_strm1_data_valid  ;

  input                                         std__mgr13__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane4_strm0_data        ;
  output                                        mgr13__std__lane4_strm0_data_valid  ;

  input                                         std__mgr13__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane4_strm1_data        ;
  output                                        mgr13__std__lane4_strm1_data_valid  ;

  input                                         std__mgr13__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane5_strm0_data        ;
  output                                        mgr13__std__lane5_strm0_data_valid  ;

  input                                         std__mgr13__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane5_strm1_data        ;
  output                                        mgr13__std__lane5_strm1_data_valid  ;

  input                                         std__mgr13__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane6_strm0_data        ;
  output                                        mgr13__std__lane6_strm0_data_valid  ;

  input                                         std__mgr13__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane6_strm1_data        ;
  output                                        mgr13__std__lane6_strm1_data_valid  ;

  input                                         std__mgr13__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane7_strm0_data        ;
  output                                        mgr13__std__lane7_strm0_data_valid  ;

  input                                         std__mgr13__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane7_strm1_data        ;
  output                                        mgr13__std__lane7_strm1_data_valid  ;

  input                                         std__mgr13__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane8_strm0_data        ;
  output                                        mgr13__std__lane8_strm0_data_valid  ;

  input                                         std__mgr13__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane8_strm1_data        ;
  output                                        mgr13__std__lane8_strm1_data_valid  ;

  input                                         std__mgr13__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane9_strm0_data        ;
  output                                        mgr13__std__lane9_strm0_data_valid  ;

  input                                         std__mgr13__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane9_strm1_data        ;
  output                                        mgr13__std__lane9_strm1_data_valid  ;

  input                                         std__mgr13__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane10_strm0_data        ;
  output                                        mgr13__std__lane10_strm0_data_valid  ;

  input                                         std__mgr13__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane10_strm1_data        ;
  output                                        mgr13__std__lane10_strm1_data_valid  ;

  input                                         std__mgr13__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane11_strm0_data        ;
  output                                        mgr13__std__lane11_strm0_data_valid  ;

  input                                         std__mgr13__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane11_strm1_data        ;
  output                                        mgr13__std__lane11_strm1_data_valid  ;

  input                                         std__mgr13__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane12_strm0_data        ;
  output                                        mgr13__std__lane12_strm0_data_valid  ;

  input                                         std__mgr13__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane12_strm1_data        ;
  output                                        mgr13__std__lane12_strm1_data_valid  ;

  input                                         std__mgr13__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane13_strm0_data        ;
  output                                        mgr13__std__lane13_strm0_data_valid  ;

  input                                         std__mgr13__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane13_strm1_data        ;
  output                                        mgr13__std__lane13_strm1_data_valid  ;

  input                                         std__mgr13__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane14_strm0_data        ;
  output                                        mgr13__std__lane14_strm0_data_valid  ;

  input                                         std__mgr13__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane14_strm1_data        ;
  output                                        mgr13__std__lane14_strm1_data_valid  ;

  input                                         std__mgr13__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane15_strm0_data        ;
  output                                        mgr13__std__lane15_strm0_data_valid  ;

  input                                         std__mgr13__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane15_strm1_data        ;
  output                                        mgr13__std__lane15_strm1_data_valid  ;

  input                                         std__mgr13__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane16_strm0_data        ;
  output                                        mgr13__std__lane16_strm0_data_valid  ;

  input                                         std__mgr13__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane16_strm1_data        ;
  output                                        mgr13__std__lane16_strm1_data_valid  ;

  input                                         std__mgr13__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane17_strm0_data        ;
  output                                        mgr13__std__lane17_strm0_data_valid  ;

  input                                         std__mgr13__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane17_strm1_data        ;
  output                                        mgr13__std__lane17_strm1_data_valid  ;

  input                                         std__mgr13__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane18_strm0_data        ;
  output                                        mgr13__std__lane18_strm0_data_valid  ;

  input                                         std__mgr13__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane18_strm1_data        ;
  output                                        mgr13__std__lane18_strm1_data_valid  ;

  input                                         std__mgr13__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane19_strm0_data        ;
  output                                        mgr13__std__lane19_strm0_data_valid  ;

  input                                         std__mgr13__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane19_strm1_data        ;
  output                                        mgr13__std__lane19_strm1_data_valid  ;

  input                                         std__mgr13__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane20_strm0_data        ;
  output                                        mgr13__std__lane20_strm0_data_valid  ;

  input                                         std__mgr13__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane20_strm1_data        ;
  output                                        mgr13__std__lane20_strm1_data_valid  ;

  input                                         std__mgr13__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane21_strm0_data        ;
  output                                        mgr13__std__lane21_strm0_data_valid  ;

  input                                         std__mgr13__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane21_strm1_data        ;
  output                                        mgr13__std__lane21_strm1_data_valid  ;

  input                                         std__mgr13__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane22_strm0_data        ;
  output                                        mgr13__std__lane22_strm0_data_valid  ;

  input                                         std__mgr13__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane22_strm1_data        ;
  output                                        mgr13__std__lane22_strm1_data_valid  ;

  input                                         std__mgr13__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane23_strm0_data        ;
  output                                        mgr13__std__lane23_strm0_data_valid  ;

  input                                         std__mgr13__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane23_strm1_data        ;
  output                                        mgr13__std__lane23_strm1_data_valid  ;

  input                                         std__mgr13__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane24_strm0_data        ;
  output                                        mgr13__std__lane24_strm0_data_valid  ;

  input                                         std__mgr13__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane24_strm1_data        ;
  output                                        mgr13__std__lane24_strm1_data_valid  ;

  input                                         std__mgr13__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane25_strm0_data        ;
  output                                        mgr13__std__lane25_strm0_data_valid  ;

  input                                         std__mgr13__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane25_strm1_data        ;
  output                                        mgr13__std__lane25_strm1_data_valid  ;

  input                                         std__mgr13__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane26_strm0_data        ;
  output                                        mgr13__std__lane26_strm0_data_valid  ;

  input                                         std__mgr13__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane26_strm1_data        ;
  output                                        mgr13__std__lane26_strm1_data_valid  ;

  input                                         std__mgr13__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane27_strm0_data        ;
  output                                        mgr13__std__lane27_strm0_data_valid  ;

  input                                         std__mgr13__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane27_strm1_data        ;
  output                                        mgr13__std__lane27_strm1_data_valid  ;

  input                                         std__mgr13__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane28_strm0_data        ;
  output                                        mgr13__std__lane28_strm0_data_valid  ;

  input                                         std__mgr13__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane28_strm1_data        ;
  output                                        mgr13__std__lane28_strm1_data_valid  ;

  input                                         std__mgr13__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane29_strm0_data        ;
  output                                        mgr13__std__lane29_strm0_data_valid  ;

  input                                         std__mgr13__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane29_strm1_data        ;
  output                                        mgr13__std__lane29_strm1_data_valid  ;

  input                                         std__mgr13__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane30_strm0_data        ;
  output                                        mgr13__std__lane30_strm0_data_valid  ;

  input                                         std__mgr13__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane30_strm1_data        ;
  output                                        mgr13__std__lane30_strm1_data_valid  ;

  input                                         std__mgr13__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane31_strm0_data        ;
  output                                        mgr13__std__lane31_strm0_data_valid  ;

  input                                         std__mgr13__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane31_strm1_data        ;
  output                                        mgr13__std__lane31_strm1_data_valid  ;

  input                                         std__mgr14__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane0_strm0_data        ;
  output                                        mgr14__std__lane0_strm0_data_valid  ;

  input                                         std__mgr14__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane0_strm1_data        ;
  output                                        mgr14__std__lane0_strm1_data_valid  ;

  input                                         std__mgr14__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane1_strm0_data        ;
  output                                        mgr14__std__lane1_strm0_data_valid  ;

  input                                         std__mgr14__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane1_strm1_data        ;
  output                                        mgr14__std__lane1_strm1_data_valid  ;

  input                                         std__mgr14__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane2_strm0_data        ;
  output                                        mgr14__std__lane2_strm0_data_valid  ;

  input                                         std__mgr14__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane2_strm1_data        ;
  output                                        mgr14__std__lane2_strm1_data_valid  ;

  input                                         std__mgr14__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane3_strm0_data        ;
  output                                        mgr14__std__lane3_strm0_data_valid  ;

  input                                         std__mgr14__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane3_strm1_data        ;
  output                                        mgr14__std__lane3_strm1_data_valid  ;

  input                                         std__mgr14__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane4_strm0_data        ;
  output                                        mgr14__std__lane4_strm0_data_valid  ;

  input                                         std__mgr14__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane4_strm1_data        ;
  output                                        mgr14__std__lane4_strm1_data_valid  ;

  input                                         std__mgr14__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane5_strm0_data        ;
  output                                        mgr14__std__lane5_strm0_data_valid  ;

  input                                         std__mgr14__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane5_strm1_data        ;
  output                                        mgr14__std__lane5_strm1_data_valid  ;

  input                                         std__mgr14__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane6_strm0_data        ;
  output                                        mgr14__std__lane6_strm0_data_valid  ;

  input                                         std__mgr14__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane6_strm1_data        ;
  output                                        mgr14__std__lane6_strm1_data_valid  ;

  input                                         std__mgr14__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane7_strm0_data        ;
  output                                        mgr14__std__lane7_strm0_data_valid  ;

  input                                         std__mgr14__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane7_strm1_data        ;
  output                                        mgr14__std__lane7_strm1_data_valid  ;

  input                                         std__mgr14__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane8_strm0_data        ;
  output                                        mgr14__std__lane8_strm0_data_valid  ;

  input                                         std__mgr14__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane8_strm1_data        ;
  output                                        mgr14__std__lane8_strm1_data_valid  ;

  input                                         std__mgr14__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane9_strm0_data        ;
  output                                        mgr14__std__lane9_strm0_data_valid  ;

  input                                         std__mgr14__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane9_strm1_data        ;
  output                                        mgr14__std__lane9_strm1_data_valid  ;

  input                                         std__mgr14__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane10_strm0_data        ;
  output                                        mgr14__std__lane10_strm0_data_valid  ;

  input                                         std__mgr14__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane10_strm1_data        ;
  output                                        mgr14__std__lane10_strm1_data_valid  ;

  input                                         std__mgr14__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane11_strm0_data        ;
  output                                        mgr14__std__lane11_strm0_data_valid  ;

  input                                         std__mgr14__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane11_strm1_data        ;
  output                                        mgr14__std__lane11_strm1_data_valid  ;

  input                                         std__mgr14__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane12_strm0_data        ;
  output                                        mgr14__std__lane12_strm0_data_valid  ;

  input                                         std__mgr14__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane12_strm1_data        ;
  output                                        mgr14__std__lane12_strm1_data_valid  ;

  input                                         std__mgr14__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane13_strm0_data        ;
  output                                        mgr14__std__lane13_strm0_data_valid  ;

  input                                         std__mgr14__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane13_strm1_data        ;
  output                                        mgr14__std__lane13_strm1_data_valid  ;

  input                                         std__mgr14__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane14_strm0_data        ;
  output                                        mgr14__std__lane14_strm0_data_valid  ;

  input                                         std__mgr14__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane14_strm1_data        ;
  output                                        mgr14__std__lane14_strm1_data_valid  ;

  input                                         std__mgr14__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane15_strm0_data        ;
  output                                        mgr14__std__lane15_strm0_data_valid  ;

  input                                         std__mgr14__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane15_strm1_data        ;
  output                                        mgr14__std__lane15_strm1_data_valid  ;

  input                                         std__mgr14__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane16_strm0_data        ;
  output                                        mgr14__std__lane16_strm0_data_valid  ;

  input                                         std__mgr14__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane16_strm1_data        ;
  output                                        mgr14__std__lane16_strm1_data_valid  ;

  input                                         std__mgr14__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane17_strm0_data        ;
  output                                        mgr14__std__lane17_strm0_data_valid  ;

  input                                         std__mgr14__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane17_strm1_data        ;
  output                                        mgr14__std__lane17_strm1_data_valid  ;

  input                                         std__mgr14__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane18_strm0_data        ;
  output                                        mgr14__std__lane18_strm0_data_valid  ;

  input                                         std__mgr14__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane18_strm1_data        ;
  output                                        mgr14__std__lane18_strm1_data_valid  ;

  input                                         std__mgr14__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane19_strm0_data        ;
  output                                        mgr14__std__lane19_strm0_data_valid  ;

  input                                         std__mgr14__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane19_strm1_data        ;
  output                                        mgr14__std__lane19_strm1_data_valid  ;

  input                                         std__mgr14__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane20_strm0_data        ;
  output                                        mgr14__std__lane20_strm0_data_valid  ;

  input                                         std__mgr14__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane20_strm1_data        ;
  output                                        mgr14__std__lane20_strm1_data_valid  ;

  input                                         std__mgr14__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane21_strm0_data        ;
  output                                        mgr14__std__lane21_strm0_data_valid  ;

  input                                         std__mgr14__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane21_strm1_data        ;
  output                                        mgr14__std__lane21_strm1_data_valid  ;

  input                                         std__mgr14__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane22_strm0_data        ;
  output                                        mgr14__std__lane22_strm0_data_valid  ;

  input                                         std__mgr14__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane22_strm1_data        ;
  output                                        mgr14__std__lane22_strm1_data_valid  ;

  input                                         std__mgr14__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane23_strm0_data        ;
  output                                        mgr14__std__lane23_strm0_data_valid  ;

  input                                         std__mgr14__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane23_strm1_data        ;
  output                                        mgr14__std__lane23_strm1_data_valid  ;

  input                                         std__mgr14__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane24_strm0_data        ;
  output                                        mgr14__std__lane24_strm0_data_valid  ;

  input                                         std__mgr14__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane24_strm1_data        ;
  output                                        mgr14__std__lane24_strm1_data_valid  ;

  input                                         std__mgr14__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane25_strm0_data        ;
  output                                        mgr14__std__lane25_strm0_data_valid  ;

  input                                         std__mgr14__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane25_strm1_data        ;
  output                                        mgr14__std__lane25_strm1_data_valid  ;

  input                                         std__mgr14__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane26_strm0_data        ;
  output                                        mgr14__std__lane26_strm0_data_valid  ;

  input                                         std__mgr14__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane26_strm1_data        ;
  output                                        mgr14__std__lane26_strm1_data_valid  ;

  input                                         std__mgr14__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane27_strm0_data        ;
  output                                        mgr14__std__lane27_strm0_data_valid  ;

  input                                         std__mgr14__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane27_strm1_data        ;
  output                                        mgr14__std__lane27_strm1_data_valid  ;

  input                                         std__mgr14__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane28_strm0_data        ;
  output                                        mgr14__std__lane28_strm0_data_valid  ;

  input                                         std__mgr14__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane28_strm1_data        ;
  output                                        mgr14__std__lane28_strm1_data_valid  ;

  input                                         std__mgr14__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane29_strm0_data        ;
  output                                        mgr14__std__lane29_strm0_data_valid  ;

  input                                         std__mgr14__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane29_strm1_data        ;
  output                                        mgr14__std__lane29_strm1_data_valid  ;

  input                                         std__mgr14__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane30_strm0_data        ;
  output                                        mgr14__std__lane30_strm0_data_valid  ;

  input                                         std__mgr14__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane30_strm1_data        ;
  output                                        mgr14__std__lane30_strm1_data_valid  ;

  input                                         std__mgr14__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane31_strm0_data        ;
  output                                        mgr14__std__lane31_strm0_data_valid  ;

  input                                         std__mgr14__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane31_strm1_data        ;
  output                                        mgr14__std__lane31_strm1_data_valid  ;

  input                                         std__mgr15__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane0_strm0_data        ;
  output                                        mgr15__std__lane0_strm0_data_valid  ;

  input                                         std__mgr15__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane0_strm1_data        ;
  output                                        mgr15__std__lane0_strm1_data_valid  ;

  input                                         std__mgr15__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane1_strm0_data        ;
  output                                        mgr15__std__lane1_strm0_data_valid  ;

  input                                         std__mgr15__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane1_strm1_data        ;
  output                                        mgr15__std__lane1_strm1_data_valid  ;

  input                                         std__mgr15__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane2_strm0_data        ;
  output                                        mgr15__std__lane2_strm0_data_valid  ;

  input                                         std__mgr15__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane2_strm1_data        ;
  output                                        mgr15__std__lane2_strm1_data_valid  ;

  input                                         std__mgr15__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane3_strm0_data        ;
  output                                        mgr15__std__lane3_strm0_data_valid  ;

  input                                         std__mgr15__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane3_strm1_data        ;
  output                                        mgr15__std__lane3_strm1_data_valid  ;

  input                                         std__mgr15__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane4_strm0_data        ;
  output                                        mgr15__std__lane4_strm0_data_valid  ;

  input                                         std__mgr15__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane4_strm1_data        ;
  output                                        mgr15__std__lane4_strm1_data_valid  ;

  input                                         std__mgr15__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane5_strm0_data        ;
  output                                        mgr15__std__lane5_strm0_data_valid  ;

  input                                         std__mgr15__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane5_strm1_data        ;
  output                                        mgr15__std__lane5_strm1_data_valid  ;

  input                                         std__mgr15__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane6_strm0_data        ;
  output                                        mgr15__std__lane6_strm0_data_valid  ;

  input                                         std__mgr15__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane6_strm1_data        ;
  output                                        mgr15__std__lane6_strm1_data_valid  ;

  input                                         std__mgr15__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane7_strm0_data        ;
  output                                        mgr15__std__lane7_strm0_data_valid  ;

  input                                         std__mgr15__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane7_strm1_data        ;
  output                                        mgr15__std__lane7_strm1_data_valid  ;

  input                                         std__mgr15__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane8_strm0_data        ;
  output                                        mgr15__std__lane8_strm0_data_valid  ;

  input                                         std__mgr15__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane8_strm1_data        ;
  output                                        mgr15__std__lane8_strm1_data_valid  ;

  input                                         std__mgr15__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane9_strm0_data        ;
  output                                        mgr15__std__lane9_strm0_data_valid  ;

  input                                         std__mgr15__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane9_strm1_data        ;
  output                                        mgr15__std__lane9_strm1_data_valid  ;

  input                                         std__mgr15__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane10_strm0_data        ;
  output                                        mgr15__std__lane10_strm0_data_valid  ;

  input                                         std__mgr15__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane10_strm1_data        ;
  output                                        mgr15__std__lane10_strm1_data_valid  ;

  input                                         std__mgr15__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane11_strm0_data        ;
  output                                        mgr15__std__lane11_strm0_data_valid  ;

  input                                         std__mgr15__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane11_strm1_data        ;
  output                                        mgr15__std__lane11_strm1_data_valid  ;

  input                                         std__mgr15__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane12_strm0_data        ;
  output                                        mgr15__std__lane12_strm0_data_valid  ;

  input                                         std__mgr15__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane12_strm1_data        ;
  output                                        mgr15__std__lane12_strm1_data_valid  ;

  input                                         std__mgr15__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane13_strm0_data        ;
  output                                        mgr15__std__lane13_strm0_data_valid  ;

  input                                         std__mgr15__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane13_strm1_data        ;
  output                                        mgr15__std__lane13_strm1_data_valid  ;

  input                                         std__mgr15__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane14_strm0_data        ;
  output                                        mgr15__std__lane14_strm0_data_valid  ;

  input                                         std__mgr15__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane14_strm1_data        ;
  output                                        mgr15__std__lane14_strm1_data_valid  ;

  input                                         std__mgr15__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane15_strm0_data        ;
  output                                        mgr15__std__lane15_strm0_data_valid  ;

  input                                         std__mgr15__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane15_strm1_data        ;
  output                                        mgr15__std__lane15_strm1_data_valid  ;

  input                                         std__mgr15__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane16_strm0_data        ;
  output                                        mgr15__std__lane16_strm0_data_valid  ;

  input                                         std__mgr15__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane16_strm1_data        ;
  output                                        mgr15__std__lane16_strm1_data_valid  ;

  input                                         std__mgr15__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane17_strm0_data        ;
  output                                        mgr15__std__lane17_strm0_data_valid  ;

  input                                         std__mgr15__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane17_strm1_data        ;
  output                                        mgr15__std__lane17_strm1_data_valid  ;

  input                                         std__mgr15__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane18_strm0_data        ;
  output                                        mgr15__std__lane18_strm0_data_valid  ;

  input                                         std__mgr15__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane18_strm1_data        ;
  output                                        mgr15__std__lane18_strm1_data_valid  ;

  input                                         std__mgr15__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane19_strm0_data        ;
  output                                        mgr15__std__lane19_strm0_data_valid  ;

  input                                         std__mgr15__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane19_strm1_data        ;
  output                                        mgr15__std__lane19_strm1_data_valid  ;

  input                                         std__mgr15__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane20_strm0_data        ;
  output                                        mgr15__std__lane20_strm0_data_valid  ;

  input                                         std__mgr15__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane20_strm1_data        ;
  output                                        mgr15__std__lane20_strm1_data_valid  ;

  input                                         std__mgr15__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane21_strm0_data        ;
  output                                        mgr15__std__lane21_strm0_data_valid  ;

  input                                         std__mgr15__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane21_strm1_data        ;
  output                                        mgr15__std__lane21_strm1_data_valid  ;

  input                                         std__mgr15__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane22_strm0_data        ;
  output                                        mgr15__std__lane22_strm0_data_valid  ;

  input                                         std__mgr15__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane22_strm1_data        ;
  output                                        mgr15__std__lane22_strm1_data_valid  ;

  input                                         std__mgr15__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane23_strm0_data        ;
  output                                        mgr15__std__lane23_strm0_data_valid  ;

  input                                         std__mgr15__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane23_strm1_data        ;
  output                                        mgr15__std__lane23_strm1_data_valid  ;

  input                                         std__mgr15__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane24_strm0_data        ;
  output                                        mgr15__std__lane24_strm0_data_valid  ;

  input                                         std__mgr15__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane24_strm1_data        ;
  output                                        mgr15__std__lane24_strm1_data_valid  ;

  input                                         std__mgr15__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane25_strm0_data        ;
  output                                        mgr15__std__lane25_strm0_data_valid  ;

  input                                         std__mgr15__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane25_strm1_data        ;
  output                                        mgr15__std__lane25_strm1_data_valid  ;

  input                                         std__mgr15__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane26_strm0_data        ;
  output                                        mgr15__std__lane26_strm0_data_valid  ;

  input                                         std__mgr15__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane26_strm1_data        ;
  output                                        mgr15__std__lane26_strm1_data_valid  ;

  input                                         std__mgr15__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane27_strm0_data        ;
  output                                        mgr15__std__lane27_strm0_data_valid  ;

  input                                         std__mgr15__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane27_strm1_data        ;
  output                                        mgr15__std__lane27_strm1_data_valid  ;

  input                                         std__mgr15__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane28_strm0_data        ;
  output                                        mgr15__std__lane28_strm0_data_valid  ;

  input                                         std__mgr15__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane28_strm1_data        ;
  output                                        mgr15__std__lane28_strm1_data_valid  ;

  input                                         std__mgr15__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane29_strm0_data        ;
  output                                        mgr15__std__lane29_strm0_data_valid  ;

  input                                         std__mgr15__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane29_strm1_data        ;
  output                                        mgr15__std__lane29_strm1_data_valid  ;

  input                                         std__mgr15__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane30_strm0_data        ;
  output                                        mgr15__std__lane30_strm0_data_valid  ;

  input                                         std__mgr15__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane30_strm1_data        ;
  output                                        mgr15__std__lane30_strm1_data_valid  ;

  input                                         std__mgr15__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane31_strm0_data        ;
  output                                        mgr15__std__lane31_strm0_data_valid  ;

  input                                         std__mgr15__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane31_strm1_data        ;
  output                                        mgr15__std__lane31_strm1_data_valid  ;

  input                                         std__mgr16__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane0_strm0_data        ;
  output                                        mgr16__std__lane0_strm0_data_valid  ;

  input                                         std__mgr16__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane0_strm1_data        ;
  output                                        mgr16__std__lane0_strm1_data_valid  ;

  input                                         std__mgr16__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane1_strm0_data        ;
  output                                        mgr16__std__lane1_strm0_data_valid  ;

  input                                         std__mgr16__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane1_strm1_data        ;
  output                                        mgr16__std__lane1_strm1_data_valid  ;

  input                                         std__mgr16__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane2_strm0_data        ;
  output                                        mgr16__std__lane2_strm0_data_valid  ;

  input                                         std__mgr16__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane2_strm1_data        ;
  output                                        mgr16__std__lane2_strm1_data_valid  ;

  input                                         std__mgr16__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane3_strm0_data        ;
  output                                        mgr16__std__lane3_strm0_data_valid  ;

  input                                         std__mgr16__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane3_strm1_data        ;
  output                                        mgr16__std__lane3_strm1_data_valid  ;

  input                                         std__mgr16__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane4_strm0_data        ;
  output                                        mgr16__std__lane4_strm0_data_valid  ;

  input                                         std__mgr16__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane4_strm1_data        ;
  output                                        mgr16__std__lane4_strm1_data_valid  ;

  input                                         std__mgr16__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane5_strm0_data        ;
  output                                        mgr16__std__lane5_strm0_data_valid  ;

  input                                         std__mgr16__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane5_strm1_data        ;
  output                                        mgr16__std__lane5_strm1_data_valid  ;

  input                                         std__mgr16__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane6_strm0_data        ;
  output                                        mgr16__std__lane6_strm0_data_valid  ;

  input                                         std__mgr16__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane6_strm1_data        ;
  output                                        mgr16__std__lane6_strm1_data_valid  ;

  input                                         std__mgr16__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane7_strm0_data        ;
  output                                        mgr16__std__lane7_strm0_data_valid  ;

  input                                         std__mgr16__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane7_strm1_data        ;
  output                                        mgr16__std__lane7_strm1_data_valid  ;

  input                                         std__mgr16__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane8_strm0_data        ;
  output                                        mgr16__std__lane8_strm0_data_valid  ;

  input                                         std__mgr16__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane8_strm1_data        ;
  output                                        mgr16__std__lane8_strm1_data_valid  ;

  input                                         std__mgr16__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane9_strm0_data        ;
  output                                        mgr16__std__lane9_strm0_data_valid  ;

  input                                         std__mgr16__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane9_strm1_data        ;
  output                                        mgr16__std__lane9_strm1_data_valid  ;

  input                                         std__mgr16__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane10_strm0_data        ;
  output                                        mgr16__std__lane10_strm0_data_valid  ;

  input                                         std__mgr16__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane10_strm1_data        ;
  output                                        mgr16__std__lane10_strm1_data_valid  ;

  input                                         std__mgr16__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane11_strm0_data        ;
  output                                        mgr16__std__lane11_strm0_data_valid  ;

  input                                         std__mgr16__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane11_strm1_data        ;
  output                                        mgr16__std__lane11_strm1_data_valid  ;

  input                                         std__mgr16__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane12_strm0_data        ;
  output                                        mgr16__std__lane12_strm0_data_valid  ;

  input                                         std__mgr16__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane12_strm1_data        ;
  output                                        mgr16__std__lane12_strm1_data_valid  ;

  input                                         std__mgr16__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane13_strm0_data        ;
  output                                        mgr16__std__lane13_strm0_data_valid  ;

  input                                         std__mgr16__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane13_strm1_data        ;
  output                                        mgr16__std__lane13_strm1_data_valid  ;

  input                                         std__mgr16__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane14_strm0_data        ;
  output                                        mgr16__std__lane14_strm0_data_valid  ;

  input                                         std__mgr16__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane14_strm1_data        ;
  output                                        mgr16__std__lane14_strm1_data_valid  ;

  input                                         std__mgr16__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane15_strm0_data        ;
  output                                        mgr16__std__lane15_strm0_data_valid  ;

  input                                         std__mgr16__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane15_strm1_data        ;
  output                                        mgr16__std__lane15_strm1_data_valid  ;

  input                                         std__mgr16__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane16_strm0_data        ;
  output                                        mgr16__std__lane16_strm0_data_valid  ;

  input                                         std__mgr16__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane16_strm1_data        ;
  output                                        mgr16__std__lane16_strm1_data_valid  ;

  input                                         std__mgr16__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane17_strm0_data        ;
  output                                        mgr16__std__lane17_strm0_data_valid  ;

  input                                         std__mgr16__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane17_strm1_data        ;
  output                                        mgr16__std__lane17_strm1_data_valid  ;

  input                                         std__mgr16__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane18_strm0_data        ;
  output                                        mgr16__std__lane18_strm0_data_valid  ;

  input                                         std__mgr16__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane18_strm1_data        ;
  output                                        mgr16__std__lane18_strm1_data_valid  ;

  input                                         std__mgr16__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane19_strm0_data        ;
  output                                        mgr16__std__lane19_strm0_data_valid  ;

  input                                         std__mgr16__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane19_strm1_data        ;
  output                                        mgr16__std__lane19_strm1_data_valid  ;

  input                                         std__mgr16__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane20_strm0_data        ;
  output                                        mgr16__std__lane20_strm0_data_valid  ;

  input                                         std__mgr16__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane20_strm1_data        ;
  output                                        mgr16__std__lane20_strm1_data_valid  ;

  input                                         std__mgr16__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane21_strm0_data        ;
  output                                        mgr16__std__lane21_strm0_data_valid  ;

  input                                         std__mgr16__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane21_strm1_data        ;
  output                                        mgr16__std__lane21_strm1_data_valid  ;

  input                                         std__mgr16__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane22_strm0_data        ;
  output                                        mgr16__std__lane22_strm0_data_valid  ;

  input                                         std__mgr16__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane22_strm1_data        ;
  output                                        mgr16__std__lane22_strm1_data_valid  ;

  input                                         std__mgr16__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane23_strm0_data        ;
  output                                        mgr16__std__lane23_strm0_data_valid  ;

  input                                         std__mgr16__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane23_strm1_data        ;
  output                                        mgr16__std__lane23_strm1_data_valid  ;

  input                                         std__mgr16__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane24_strm0_data        ;
  output                                        mgr16__std__lane24_strm0_data_valid  ;

  input                                         std__mgr16__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane24_strm1_data        ;
  output                                        mgr16__std__lane24_strm1_data_valid  ;

  input                                         std__mgr16__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane25_strm0_data        ;
  output                                        mgr16__std__lane25_strm0_data_valid  ;

  input                                         std__mgr16__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane25_strm1_data        ;
  output                                        mgr16__std__lane25_strm1_data_valid  ;

  input                                         std__mgr16__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane26_strm0_data        ;
  output                                        mgr16__std__lane26_strm0_data_valid  ;

  input                                         std__mgr16__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane26_strm1_data        ;
  output                                        mgr16__std__lane26_strm1_data_valid  ;

  input                                         std__mgr16__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane27_strm0_data        ;
  output                                        mgr16__std__lane27_strm0_data_valid  ;

  input                                         std__mgr16__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane27_strm1_data        ;
  output                                        mgr16__std__lane27_strm1_data_valid  ;

  input                                         std__mgr16__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane28_strm0_data        ;
  output                                        mgr16__std__lane28_strm0_data_valid  ;

  input                                         std__mgr16__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane28_strm1_data        ;
  output                                        mgr16__std__lane28_strm1_data_valid  ;

  input                                         std__mgr16__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane29_strm0_data        ;
  output                                        mgr16__std__lane29_strm0_data_valid  ;

  input                                         std__mgr16__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane29_strm1_data        ;
  output                                        mgr16__std__lane29_strm1_data_valid  ;

  input                                         std__mgr16__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane30_strm0_data        ;
  output                                        mgr16__std__lane30_strm0_data_valid  ;

  input                                         std__mgr16__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane30_strm1_data        ;
  output                                        mgr16__std__lane30_strm1_data_valid  ;

  input                                         std__mgr16__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane31_strm0_data        ;
  output                                        mgr16__std__lane31_strm0_data_valid  ;

  input                                         std__mgr16__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane31_strm1_data        ;
  output                                        mgr16__std__lane31_strm1_data_valid  ;

  input                                         std__mgr17__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane0_strm0_data        ;
  output                                        mgr17__std__lane0_strm0_data_valid  ;

  input                                         std__mgr17__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane0_strm1_data        ;
  output                                        mgr17__std__lane0_strm1_data_valid  ;

  input                                         std__mgr17__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane1_strm0_data        ;
  output                                        mgr17__std__lane1_strm0_data_valid  ;

  input                                         std__mgr17__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane1_strm1_data        ;
  output                                        mgr17__std__lane1_strm1_data_valid  ;

  input                                         std__mgr17__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane2_strm0_data        ;
  output                                        mgr17__std__lane2_strm0_data_valid  ;

  input                                         std__mgr17__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane2_strm1_data        ;
  output                                        mgr17__std__lane2_strm1_data_valid  ;

  input                                         std__mgr17__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane3_strm0_data        ;
  output                                        mgr17__std__lane3_strm0_data_valid  ;

  input                                         std__mgr17__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane3_strm1_data        ;
  output                                        mgr17__std__lane3_strm1_data_valid  ;

  input                                         std__mgr17__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane4_strm0_data        ;
  output                                        mgr17__std__lane4_strm0_data_valid  ;

  input                                         std__mgr17__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane4_strm1_data        ;
  output                                        mgr17__std__lane4_strm1_data_valid  ;

  input                                         std__mgr17__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane5_strm0_data        ;
  output                                        mgr17__std__lane5_strm0_data_valid  ;

  input                                         std__mgr17__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane5_strm1_data        ;
  output                                        mgr17__std__lane5_strm1_data_valid  ;

  input                                         std__mgr17__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane6_strm0_data        ;
  output                                        mgr17__std__lane6_strm0_data_valid  ;

  input                                         std__mgr17__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane6_strm1_data        ;
  output                                        mgr17__std__lane6_strm1_data_valid  ;

  input                                         std__mgr17__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane7_strm0_data        ;
  output                                        mgr17__std__lane7_strm0_data_valid  ;

  input                                         std__mgr17__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane7_strm1_data        ;
  output                                        mgr17__std__lane7_strm1_data_valid  ;

  input                                         std__mgr17__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane8_strm0_data        ;
  output                                        mgr17__std__lane8_strm0_data_valid  ;

  input                                         std__mgr17__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane8_strm1_data        ;
  output                                        mgr17__std__lane8_strm1_data_valid  ;

  input                                         std__mgr17__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane9_strm0_data        ;
  output                                        mgr17__std__lane9_strm0_data_valid  ;

  input                                         std__mgr17__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane9_strm1_data        ;
  output                                        mgr17__std__lane9_strm1_data_valid  ;

  input                                         std__mgr17__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane10_strm0_data        ;
  output                                        mgr17__std__lane10_strm0_data_valid  ;

  input                                         std__mgr17__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane10_strm1_data        ;
  output                                        mgr17__std__lane10_strm1_data_valid  ;

  input                                         std__mgr17__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane11_strm0_data        ;
  output                                        mgr17__std__lane11_strm0_data_valid  ;

  input                                         std__mgr17__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane11_strm1_data        ;
  output                                        mgr17__std__lane11_strm1_data_valid  ;

  input                                         std__mgr17__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane12_strm0_data        ;
  output                                        mgr17__std__lane12_strm0_data_valid  ;

  input                                         std__mgr17__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane12_strm1_data        ;
  output                                        mgr17__std__lane12_strm1_data_valid  ;

  input                                         std__mgr17__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane13_strm0_data        ;
  output                                        mgr17__std__lane13_strm0_data_valid  ;

  input                                         std__mgr17__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane13_strm1_data        ;
  output                                        mgr17__std__lane13_strm1_data_valid  ;

  input                                         std__mgr17__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane14_strm0_data        ;
  output                                        mgr17__std__lane14_strm0_data_valid  ;

  input                                         std__mgr17__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane14_strm1_data        ;
  output                                        mgr17__std__lane14_strm1_data_valid  ;

  input                                         std__mgr17__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane15_strm0_data        ;
  output                                        mgr17__std__lane15_strm0_data_valid  ;

  input                                         std__mgr17__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane15_strm1_data        ;
  output                                        mgr17__std__lane15_strm1_data_valid  ;

  input                                         std__mgr17__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane16_strm0_data        ;
  output                                        mgr17__std__lane16_strm0_data_valid  ;

  input                                         std__mgr17__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane16_strm1_data        ;
  output                                        mgr17__std__lane16_strm1_data_valid  ;

  input                                         std__mgr17__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane17_strm0_data        ;
  output                                        mgr17__std__lane17_strm0_data_valid  ;

  input                                         std__mgr17__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane17_strm1_data        ;
  output                                        mgr17__std__lane17_strm1_data_valid  ;

  input                                         std__mgr17__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane18_strm0_data        ;
  output                                        mgr17__std__lane18_strm0_data_valid  ;

  input                                         std__mgr17__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane18_strm1_data        ;
  output                                        mgr17__std__lane18_strm1_data_valid  ;

  input                                         std__mgr17__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane19_strm0_data        ;
  output                                        mgr17__std__lane19_strm0_data_valid  ;

  input                                         std__mgr17__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane19_strm1_data        ;
  output                                        mgr17__std__lane19_strm1_data_valid  ;

  input                                         std__mgr17__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane20_strm0_data        ;
  output                                        mgr17__std__lane20_strm0_data_valid  ;

  input                                         std__mgr17__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane20_strm1_data        ;
  output                                        mgr17__std__lane20_strm1_data_valid  ;

  input                                         std__mgr17__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane21_strm0_data        ;
  output                                        mgr17__std__lane21_strm0_data_valid  ;

  input                                         std__mgr17__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane21_strm1_data        ;
  output                                        mgr17__std__lane21_strm1_data_valid  ;

  input                                         std__mgr17__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane22_strm0_data        ;
  output                                        mgr17__std__lane22_strm0_data_valid  ;

  input                                         std__mgr17__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane22_strm1_data        ;
  output                                        mgr17__std__lane22_strm1_data_valid  ;

  input                                         std__mgr17__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane23_strm0_data        ;
  output                                        mgr17__std__lane23_strm0_data_valid  ;

  input                                         std__mgr17__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane23_strm1_data        ;
  output                                        mgr17__std__lane23_strm1_data_valid  ;

  input                                         std__mgr17__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane24_strm0_data        ;
  output                                        mgr17__std__lane24_strm0_data_valid  ;

  input                                         std__mgr17__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane24_strm1_data        ;
  output                                        mgr17__std__lane24_strm1_data_valid  ;

  input                                         std__mgr17__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane25_strm0_data        ;
  output                                        mgr17__std__lane25_strm0_data_valid  ;

  input                                         std__mgr17__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane25_strm1_data        ;
  output                                        mgr17__std__lane25_strm1_data_valid  ;

  input                                         std__mgr17__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane26_strm0_data        ;
  output                                        mgr17__std__lane26_strm0_data_valid  ;

  input                                         std__mgr17__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane26_strm1_data        ;
  output                                        mgr17__std__lane26_strm1_data_valid  ;

  input                                         std__mgr17__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane27_strm0_data        ;
  output                                        mgr17__std__lane27_strm0_data_valid  ;

  input                                         std__mgr17__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane27_strm1_data        ;
  output                                        mgr17__std__lane27_strm1_data_valid  ;

  input                                         std__mgr17__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane28_strm0_data        ;
  output                                        mgr17__std__lane28_strm0_data_valid  ;

  input                                         std__mgr17__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane28_strm1_data        ;
  output                                        mgr17__std__lane28_strm1_data_valid  ;

  input                                         std__mgr17__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane29_strm0_data        ;
  output                                        mgr17__std__lane29_strm0_data_valid  ;

  input                                         std__mgr17__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane29_strm1_data        ;
  output                                        mgr17__std__lane29_strm1_data_valid  ;

  input                                         std__mgr17__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane30_strm0_data        ;
  output                                        mgr17__std__lane30_strm0_data_valid  ;

  input                                         std__mgr17__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane30_strm1_data        ;
  output                                        mgr17__std__lane30_strm1_data_valid  ;

  input                                         std__mgr17__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane31_strm0_data        ;
  output                                        mgr17__std__lane31_strm0_data_valid  ;

  input                                         std__mgr17__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane31_strm1_data        ;
  output                                        mgr17__std__lane31_strm1_data_valid  ;

  input                                         std__mgr18__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane0_strm0_data        ;
  output                                        mgr18__std__lane0_strm0_data_valid  ;

  input                                         std__mgr18__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane0_strm1_data        ;
  output                                        mgr18__std__lane0_strm1_data_valid  ;

  input                                         std__mgr18__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane1_strm0_data        ;
  output                                        mgr18__std__lane1_strm0_data_valid  ;

  input                                         std__mgr18__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane1_strm1_data        ;
  output                                        mgr18__std__lane1_strm1_data_valid  ;

  input                                         std__mgr18__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane2_strm0_data        ;
  output                                        mgr18__std__lane2_strm0_data_valid  ;

  input                                         std__mgr18__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane2_strm1_data        ;
  output                                        mgr18__std__lane2_strm1_data_valid  ;

  input                                         std__mgr18__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane3_strm0_data        ;
  output                                        mgr18__std__lane3_strm0_data_valid  ;

  input                                         std__mgr18__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane3_strm1_data        ;
  output                                        mgr18__std__lane3_strm1_data_valid  ;

  input                                         std__mgr18__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane4_strm0_data        ;
  output                                        mgr18__std__lane4_strm0_data_valid  ;

  input                                         std__mgr18__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane4_strm1_data        ;
  output                                        mgr18__std__lane4_strm1_data_valid  ;

  input                                         std__mgr18__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane5_strm0_data        ;
  output                                        mgr18__std__lane5_strm0_data_valid  ;

  input                                         std__mgr18__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane5_strm1_data        ;
  output                                        mgr18__std__lane5_strm1_data_valid  ;

  input                                         std__mgr18__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane6_strm0_data        ;
  output                                        mgr18__std__lane6_strm0_data_valid  ;

  input                                         std__mgr18__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane6_strm1_data        ;
  output                                        mgr18__std__lane6_strm1_data_valid  ;

  input                                         std__mgr18__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane7_strm0_data        ;
  output                                        mgr18__std__lane7_strm0_data_valid  ;

  input                                         std__mgr18__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane7_strm1_data        ;
  output                                        mgr18__std__lane7_strm1_data_valid  ;

  input                                         std__mgr18__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane8_strm0_data        ;
  output                                        mgr18__std__lane8_strm0_data_valid  ;

  input                                         std__mgr18__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane8_strm1_data        ;
  output                                        mgr18__std__lane8_strm1_data_valid  ;

  input                                         std__mgr18__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane9_strm0_data        ;
  output                                        mgr18__std__lane9_strm0_data_valid  ;

  input                                         std__mgr18__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane9_strm1_data        ;
  output                                        mgr18__std__lane9_strm1_data_valid  ;

  input                                         std__mgr18__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane10_strm0_data        ;
  output                                        mgr18__std__lane10_strm0_data_valid  ;

  input                                         std__mgr18__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane10_strm1_data        ;
  output                                        mgr18__std__lane10_strm1_data_valid  ;

  input                                         std__mgr18__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane11_strm0_data        ;
  output                                        mgr18__std__lane11_strm0_data_valid  ;

  input                                         std__mgr18__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane11_strm1_data        ;
  output                                        mgr18__std__lane11_strm1_data_valid  ;

  input                                         std__mgr18__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane12_strm0_data        ;
  output                                        mgr18__std__lane12_strm0_data_valid  ;

  input                                         std__mgr18__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane12_strm1_data        ;
  output                                        mgr18__std__lane12_strm1_data_valid  ;

  input                                         std__mgr18__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane13_strm0_data        ;
  output                                        mgr18__std__lane13_strm0_data_valid  ;

  input                                         std__mgr18__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane13_strm1_data        ;
  output                                        mgr18__std__lane13_strm1_data_valid  ;

  input                                         std__mgr18__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane14_strm0_data        ;
  output                                        mgr18__std__lane14_strm0_data_valid  ;

  input                                         std__mgr18__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane14_strm1_data        ;
  output                                        mgr18__std__lane14_strm1_data_valid  ;

  input                                         std__mgr18__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane15_strm0_data        ;
  output                                        mgr18__std__lane15_strm0_data_valid  ;

  input                                         std__mgr18__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane15_strm1_data        ;
  output                                        mgr18__std__lane15_strm1_data_valid  ;

  input                                         std__mgr18__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane16_strm0_data        ;
  output                                        mgr18__std__lane16_strm0_data_valid  ;

  input                                         std__mgr18__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane16_strm1_data        ;
  output                                        mgr18__std__lane16_strm1_data_valid  ;

  input                                         std__mgr18__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane17_strm0_data        ;
  output                                        mgr18__std__lane17_strm0_data_valid  ;

  input                                         std__mgr18__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane17_strm1_data        ;
  output                                        mgr18__std__lane17_strm1_data_valid  ;

  input                                         std__mgr18__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane18_strm0_data        ;
  output                                        mgr18__std__lane18_strm0_data_valid  ;

  input                                         std__mgr18__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane18_strm1_data        ;
  output                                        mgr18__std__lane18_strm1_data_valid  ;

  input                                         std__mgr18__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane19_strm0_data        ;
  output                                        mgr18__std__lane19_strm0_data_valid  ;

  input                                         std__mgr18__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane19_strm1_data        ;
  output                                        mgr18__std__lane19_strm1_data_valid  ;

  input                                         std__mgr18__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane20_strm0_data        ;
  output                                        mgr18__std__lane20_strm0_data_valid  ;

  input                                         std__mgr18__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane20_strm1_data        ;
  output                                        mgr18__std__lane20_strm1_data_valid  ;

  input                                         std__mgr18__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane21_strm0_data        ;
  output                                        mgr18__std__lane21_strm0_data_valid  ;

  input                                         std__mgr18__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane21_strm1_data        ;
  output                                        mgr18__std__lane21_strm1_data_valid  ;

  input                                         std__mgr18__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane22_strm0_data        ;
  output                                        mgr18__std__lane22_strm0_data_valid  ;

  input                                         std__mgr18__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane22_strm1_data        ;
  output                                        mgr18__std__lane22_strm1_data_valid  ;

  input                                         std__mgr18__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane23_strm0_data        ;
  output                                        mgr18__std__lane23_strm0_data_valid  ;

  input                                         std__mgr18__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane23_strm1_data        ;
  output                                        mgr18__std__lane23_strm1_data_valid  ;

  input                                         std__mgr18__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane24_strm0_data        ;
  output                                        mgr18__std__lane24_strm0_data_valid  ;

  input                                         std__mgr18__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane24_strm1_data        ;
  output                                        mgr18__std__lane24_strm1_data_valid  ;

  input                                         std__mgr18__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane25_strm0_data        ;
  output                                        mgr18__std__lane25_strm0_data_valid  ;

  input                                         std__mgr18__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane25_strm1_data        ;
  output                                        mgr18__std__lane25_strm1_data_valid  ;

  input                                         std__mgr18__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane26_strm0_data        ;
  output                                        mgr18__std__lane26_strm0_data_valid  ;

  input                                         std__mgr18__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane26_strm1_data        ;
  output                                        mgr18__std__lane26_strm1_data_valid  ;

  input                                         std__mgr18__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane27_strm0_data        ;
  output                                        mgr18__std__lane27_strm0_data_valid  ;

  input                                         std__mgr18__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane27_strm1_data        ;
  output                                        mgr18__std__lane27_strm1_data_valid  ;

  input                                         std__mgr18__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane28_strm0_data        ;
  output                                        mgr18__std__lane28_strm0_data_valid  ;

  input                                         std__mgr18__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane28_strm1_data        ;
  output                                        mgr18__std__lane28_strm1_data_valid  ;

  input                                         std__mgr18__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane29_strm0_data        ;
  output                                        mgr18__std__lane29_strm0_data_valid  ;

  input                                         std__mgr18__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane29_strm1_data        ;
  output                                        mgr18__std__lane29_strm1_data_valid  ;

  input                                         std__mgr18__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane30_strm0_data        ;
  output                                        mgr18__std__lane30_strm0_data_valid  ;

  input                                         std__mgr18__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane30_strm1_data        ;
  output                                        mgr18__std__lane30_strm1_data_valid  ;

  input                                         std__mgr18__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane31_strm0_data        ;
  output                                        mgr18__std__lane31_strm0_data_valid  ;

  input                                         std__mgr18__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane31_strm1_data        ;
  output                                        mgr18__std__lane31_strm1_data_valid  ;

  input                                         std__mgr19__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane0_strm0_data        ;
  output                                        mgr19__std__lane0_strm0_data_valid  ;

  input                                         std__mgr19__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane0_strm1_data        ;
  output                                        mgr19__std__lane0_strm1_data_valid  ;

  input                                         std__mgr19__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane1_strm0_data        ;
  output                                        mgr19__std__lane1_strm0_data_valid  ;

  input                                         std__mgr19__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane1_strm1_data        ;
  output                                        mgr19__std__lane1_strm1_data_valid  ;

  input                                         std__mgr19__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane2_strm0_data        ;
  output                                        mgr19__std__lane2_strm0_data_valid  ;

  input                                         std__mgr19__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane2_strm1_data        ;
  output                                        mgr19__std__lane2_strm1_data_valid  ;

  input                                         std__mgr19__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane3_strm0_data        ;
  output                                        mgr19__std__lane3_strm0_data_valid  ;

  input                                         std__mgr19__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane3_strm1_data        ;
  output                                        mgr19__std__lane3_strm1_data_valid  ;

  input                                         std__mgr19__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane4_strm0_data        ;
  output                                        mgr19__std__lane4_strm0_data_valid  ;

  input                                         std__mgr19__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane4_strm1_data        ;
  output                                        mgr19__std__lane4_strm1_data_valid  ;

  input                                         std__mgr19__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane5_strm0_data        ;
  output                                        mgr19__std__lane5_strm0_data_valid  ;

  input                                         std__mgr19__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane5_strm1_data        ;
  output                                        mgr19__std__lane5_strm1_data_valid  ;

  input                                         std__mgr19__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane6_strm0_data        ;
  output                                        mgr19__std__lane6_strm0_data_valid  ;

  input                                         std__mgr19__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane6_strm1_data        ;
  output                                        mgr19__std__lane6_strm1_data_valid  ;

  input                                         std__mgr19__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane7_strm0_data        ;
  output                                        mgr19__std__lane7_strm0_data_valid  ;

  input                                         std__mgr19__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane7_strm1_data        ;
  output                                        mgr19__std__lane7_strm1_data_valid  ;

  input                                         std__mgr19__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane8_strm0_data        ;
  output                                        mgr19__std__lane8_strm0_data_valid  ;

  input                                         std__mgr19__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane8_strm1_data        ;
  output                                        mgr19__std__lane8_strm1_data_valid  ;

  input                                         std__mgr19__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane9_strm0_data        ;
  output                                        mgr19__std__lane9_strm0_data_valid  ;

  input                                         std__mgr19__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane9_strm1_data        ;
  output                                        mgr19__std__lane9_strm1_data_valid  ;

  input                                         std__mgr19__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane10_strm0_data        ;
  output                                        mgr19__std__lane10_strm0_data_valid  ;

  input                                         std__mgr19__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane10_strm1_data        ;
  output                                        mgr19__std__lane10_strm1_data_valid  ;

  input                                         std__mgr19__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane11_strm0_data        ;
  output                                        mgr19__std__lane11_strm0_data_valid  ;

  input                                         std__mgr19__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane11_strm1_data        ;
  output                                        mgr19__std__lane11_strm1_data_valid  ;

  input                                         std__mgr19__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane12_strm0_data        ;
  output                                        mgr19__std__lane12_strm0_data_valid  ;

  input                                         std__mgr19__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane12_strm1_data        ;
  output                                        mgr19__std__lane12_strm1_data_valid  ;

  input                                         std__mgr19__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane13_strm0_data        ;
  output                                        mgr19__std__lane13_strm0_data_valid  ;

  input                                         std__mgr19__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane13_strm1_data        ;
  output                                        mgr19__std__lane13_strm1_data_valid  ;

  input                                         std__mgr19__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane14_strm0_data        ;
  output                                        mgr19__std__lane14_strm0_data_valid  ;

  input                                         std__mgr19__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane14_strm1_data        ;
  output                                        mgr19__std__lane14_strm1_data_valid  ;

  input                                         std__mgr19__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane15_strm0_data        ;
  output                                        mgr19__std__lane15_strm0_data_valid  ;

  input                                         std__mgr19__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane15_strm1_data        ;
  output                                        mgr19__std__lane15_strm1_data_valid  ;

  input                                         std__mgr19__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane16_strm0_data        ;
  output                                        mgr19__std__lane16_strm0_data_valid  ;

  input                                         std__mgr19__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane16_strm1_data        ;
  output                                        mgr19__std__lane16_strm1_data_valid  ;

  input                                         std__mgr19__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane17_strm0_data        ;
  output                                        mgr19__std__lane17_strm0_data_valid  ;

  input                                         std__mgr19__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane17_strm1_data        ;
  output                                        mgr19__std__lane17_strm1_data_valid  ;

  input                                         std__mgr19__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane18_strm0_data        ;
  output                                        mgr19__std__lane18_strm0_data_valid  ;

  input                                         std__mgr19__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane18_strm1_data        ;
  output                                        mgr19__std__lane18_strm1_data_valid  ;

  input                                         std__mgr19__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane19_strm0_data        ;
  output                                        mgr19__std__lane19_strm0_data_valid  ;

  input                                         std__mgr19__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane19_strm1_data        ;
  output                                        mgr19__std__lane19_strm1_data_valid  ;

  input                                         std__mgr19__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane20_strm0_data        ;
  output                                        mgr19__std__lane20_strm0_data_valid  ;

  input                                         std__mgr19__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane20_strm1_data        ;
  output                                        mgr19__std__lane20_strm1_data_valid  ;

  input                                         std__mgr19__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane21_strm0_data        ;
  output                                        mgr19__std__lane21_strm0_data_valid  ;

  input                                         std__mgr19__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane21_strm1_data        ;
  output                                        mgr19__std__lane21_strm1_data_valid  ;

  input                                         std__mgr19__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane22_strm0_data        ;
  output                                        mgr19__std__lane22_strm0_data_valid  ;

  input                                         std__mgr19__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane22_strm1_data        ;
  output                                        mgr19__std__lane22_strm1_data_valid  ;

  input                                         std__mgr19__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane23_strm0_data        ;
  output                                        mgr19__std__lane23_strm0_data_valid  ;

  input                                         std__mgr19__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane23_strm1_data        ;
  output                                        mgr19__std__lane23_strm1_data_valid  ;

  input                                         std__mgr19__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane24_strm0_data        ;
  output                                        mgr19__std__lane24_strm0_data_valid  ;

  input                                         std__mgr19__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane24_strm1_data        ;
  output                                        mgr19__std__lane24_strm1_data_valid  ;

  input                                         std__mgr19__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane25_strm0_data        ;
  output                                        mgr19__std__lane25_strm0_data_valid  ;

  input                                         std__mgr19__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane25_strm1_data        ;
  output                                        mgr19__std__lane25_strm1_data_valid  ;

  input                                         std__mgr19__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane26_strm0_data        ;
  output                                        mgr19__std__lane26_strm0_data_valid  ;

  input                                         std__mgr19__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane26_strm1_data        ;
  output                                        mgr19__std__lane26_strm1_data_valid  ;

  input                                         std__mgr19__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane27_strm0_data        ;
  output                                        mgr19__std__lane27_strm0_data_valid  ;

  input                                         std__mgr19__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane27_strm1_data        ;
  output                                        mgr19__std__lane27_strm1_data_valid  ;

  input                                         std__mgr19__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane28_strm0_data        ;
  output                                        mgr19__std__lane28_strm0_data_valid  ;

  input                                         std__mgr19__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane28_strm1_data        ;
  output                                        mgr19__std__lane28_strm1_data_valid  ;

  input                                         std__mgr19__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane29_strm0_data        ;
  output                                        mgr19__std__lane29_strm0_data_valid  ;

  input                                         std__mgr19__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane29_strm1_data        ;
  output                                        mgr19__std__lane29_strm1_data_valid  ;

  input                                         std__mgr19__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane30_strm0_data        ;
  output                                        mgr19__std__lane30_strm0_data_valid  ;

  input                                         std__mgr19__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane30_strm1_data        ;
  output                                        mgr19__std__lane30_strm1_data_valid  ;

  input                                         std__mgr19__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane31_strm0_data        ;
  output                                        mgr19__std__lane31_strm0_data_valid  ;

  input                                         std__mgr19__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane31_strm1_data        ;
  output                                        mgr19__std__lane31_strm1_data_valid  ;

  input                                         std__mgr20__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane0_strm0_data        ;
  output                                        mgr20__std__lane0_strm0_data_valid  ;

  input                                         std__mgr20__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane0_strm1_data        ;
  output                                        mgr20__std__lane0_strm1_data_valid  ;

  input                                         std__mgr20__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane1_strm0_data        ;
  output                                        mgr20__std__lane1_strm0_data_valid  ;

  input                                         std__mgr20__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane1_strm1_data        ;
  output                                        mgr20__std__lane1_strm1_data_valid  ;

  input                                         std__mgr20__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane2_strm0_data        ;
  output                                        mgr20__std__lane2_strm0_data_valid  ;

  input                                         std__mgr20__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane2_strm1_data        ;
  output                                        mgr20__std__lane2_strm1_data_valid  ;

  input                                         std__mgr20__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane3_strm0_data        ;
  output                                        mgr20__std__lane3_strm0_data_valid  ;

  input                                         std__mgr20__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane3_strm1_data        ;
  output                                        mgr20__std__lane3_strm1_data_valid  ;

  input                                         std__mgr20__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane4_strm0_data        ;
  output                                        mgr20__std__lane4_strm0_data_valid  ;

  input                                         std__mgr20__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane4_strm1_data        ;
  output                                        mgr20__std__lane4_strm1_data_valid  ;

  input                                         std__mgr20__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane5_strm0_data        ;
  output                                        mgr20__std__lane5_strm0_data_valid  ;

  input                                         std__mgr20__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane5_strm1_data        ;
  output                                        mgr20__std__lane5_strm1_data_valid  ;

  input                                         std__mgr20__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane6_strm0_data        ;
  output                                        mgr20__std__lane6_strm0_data_valid  ;

  input                                         std__mgr20__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane6_strm1_data        ;
  output                                        mgr20__std__lane6_strm1_data_valid  ;

  input                                         std__mgr20__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane7_strm0_data        ;
  output                                        mgr20__std__lane7_strm0_data_valid  ;

  input                                         std__mgr20__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane7_strm1_data        ;
  output                                        mgr20__std__lane7_strm1_data_valid  ;

  input                                         std__mgr20__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane8_strm0_data        ;
  output                                        mgr20__std__lane8_strm0_data_valid  ;

  input                                         std__mgr20__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane8_strm1_data        ;
  output                                        mgr20__std__lane8_strm1_data_valid  ;

  input                                         std__mgr20__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane9_strm0_data        ;
  output                                        mgr20__std__lane9_strm0_data_valid  ;

  input                                         std__mgr20__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane9_strm1_data        ;
  output                                        mgr20__std__lane9_strm1_data_valid  ;

  input                                         std__mgr20__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane10_strm0_data        ;
  output                                        mgr20__std__lane10_strm0_data_valid  ;

  input                                         std__mgr20__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane10_strm1_data        ;
  output                                        mgr20__std__lane10_strm1_data_valid  ;

  input                                         std__mgr20__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane11_strm0_data        ;
  output                                        mgr20__std__lane11_strm0_data_valid  ;

  input                                         std__mgr20__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane11_strm1_data        ;
  output                                        mgr20__std__lane11_strm1_data_valid  ;

  input                                         std__mgr20__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane12_strm0_data        ;
  output                                        mgr20__std__lane12_strm0_data_valid  ;

  input                                         std__mgr20__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane12_strm1_data        ;
  output                                        mgr20__std__lane12_strm1_data_valid  ;

  input                                         std__mgr20__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane13_strm0_data        ;
  output                                        mgr20__std__lane13_strm0_data_valid  ;

  input                                         std__mgr20__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane13_strm1_data        ;
  output                                        mgr20__std__lane13_strm1_data_valid  ;

  input                                         std__mgr20__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane14_strm0_data        ;
  output                                        mgr20__std__lane14_strm0_data_valid  ;

  input                                         std__mgr20__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane14_strm1_data        ;
  output                                        mgr20__std__lane14_strm1_data_valid  ;

  input                                         std__mgr20__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane15_strm0_data        ;
  output                                        mgr20__std__lane15_strm0_data_valid  ;

  input                                         std__mgr20__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane15_strm1_data        ;
  output                                        mgr20__std__lane15_strm1_data_valid  ;

  input                                         std__mgr20__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane16_strm0_data        ;
  output                                        mgr20__std__lane16_strm0_data_valid  ;

  input                                         std__mgr20__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane16_strm1_data        ;
  output                                        mgr20__std__lane16_strm1_data_valid  ;

  input                                         std__mgr20__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane17_strm0_data        ;
  output                                        mgr20__std__lane17_strm0_data_valid  ;

  input                                         std__mgr20__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane17_strm1_data        ;
  output                                        mgr20__std__lane17_strm1_data_valid  ;

  input                                         std__mgr20__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane18_strm0_data        ;
  output                                        mgr20__std__lane18_strm0_data_valid  ;

  input                                         std__mgr20__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane18_strm1_data        ;
  output                                        mgr20__std__lane18_strm1_data_valid  ;

  input                                         std__mgr20__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane19_strm0_data        ;
  output                                        mgr20__std__lane19_strm0_data_valid  ;

  input                                         std__mgr20__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane19_strm1_data        ;
  output                                        mgr20__std__lane19_strm1_data_valid  ;

  input                                         std__mgr20__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane20_strm0_data        ;
  output                                        mgr20__std__lane20_strm0_data_valid  ;

  input                                         std__mgr20__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane20_strm1_data        ;
  output                                        mgr20__std__lane20_strm1_data_valid  ;

  input                                         std__mgr20__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane21_strm0_data        ;
  output                                        mgr20__std__lane21_strm0_data_valid  ;

  input                                         std__mgr20__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane21_strm1_data        ;
  output                                        mgr20__std__lane21_strm1_data_valid  ;

  input                                         std__mgr20__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane22_strm0_data        ;
  output                                        mgr20__std__lane22_strm0_data_valid  ;

  input                                         std__mgr20__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane22_strm1_data        ;
  output                                        mgr20__std__lane22_strm1_data_valid  ;

  input                                         std__mgr20__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane23_strm0_data        ;
  output                                        mgr20__std__lane23_strm0_data_valid  ;

  input                                         std__mgr20__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane23_strm1_data        ;
  output                                        mgr20__std__lane23_strm1_data_valid  ;

  input                                         std__mgr20__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane24_strm0_data        ;
  output                                        mgr20__std__lane24_strm0_data_valid  ;

  input                                         std__mgr20__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane24_strm1_data        ;
  output                                        mgr20__std__lane24_strm1_data_valid  ;

  input                                         std__mgr20__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane25_strm0_data        ;
  output                                        mgr20__std__lane25_strm0_data_valid  ;

  input                                         std__mgr20__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane25_strm1_data        ;
  output                                        mgr20__std__lane25_strm1_data_valid  ;

  input                                         std__mgr20__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane26_strm0_data        ;
  output                                        mgr20__std__lane26_strm0_data_valid  ;

  input                                         std__mgr20__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane26_strm1_data        ;
  output                                        mgr20__std__lane26_strm1_data_valid  ;

  input                                         std__mgr20__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane27_strm0_data        ;
  output                                        mgr20__std__lane27_strm0_data_valid  ;

  input                                         std__mgr20__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane27_strm1_data        ;
  output                                        mgr20__std__lane27_strm1_data_valid  ;

  input                                         std__mgr20__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane28_strm0_data        ;
  output                                        mgr20__std__lane28_strm0_data_valid  ;

  input                                         std__mgr20__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane28_strm1_data        ;
  output                                        mgr20__std__lane28_strm1_data_valid  ;

  input                                         std__mgr20__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane29_strm0_data        ;
  output                                        mgr20__std__lane29_strm0_data_valid  ;

  input                                         std__mgr20__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane29_strm1_data        ;
  output                                        mgr20__std__lane29_strm1_data_valid  ;

  input                                         std__mgr20__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane30_strm0_data        ;
  output                                        mgr20__std__lane30_strm0_data_valid  ;

  input                                         std__mgr20__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane30_strm1_data        ;
  output                                        mgr20__std__lane30_strm1_data_valid  ;

  input                                         std__mgr20__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane31_strm0_data        ;
  output                                        mgr20__std__lane31_strm0_data_valid  ;

  input                                         std__mgr20__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane31_strm1_data        ;
  output                                        mgr20__std__lane31_strm1_data_valid  ;

  input                                         std__mgr21__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane0_strm0_data        ;
  output                                        mgr21__std__lane0_strm0_data_valid  ;

  input                                         std__mgr21__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane0_strm1_data        ;
  output                                        mgr21__std__lane0_strm1_data_valid  ;

  input                                         std__mgr21__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane1_strm0_data        ;
  output                                        mgr21__std__lane1_strm0_data_valid  ;

  input                                         std__mgr21__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane1_strm1_data        ;
  output                                        mgr21__std__lane1_strm1_data_valid  ;

  input                                         std__mgr21__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane2_strm0_data        ;
  output                                        mgr21__std__lane2_strm0_data_valid  ;

  input                                         std__mgr21__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane2_strm1_data        ;
  output                                        mgr21__std__lane2_strm1_data_valid  ;

  input                                         std__mgr21__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane3_strm0_data        ;
  output                                        mgr21__std__lane3_strm0_data_valid  ;

  input                                         std__mgr21__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane3_strm1_data        ;
  output                                        mgr21__std__lane3_strm1_data_valid  ;

  input                                         std__mgr21__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane4_strm0_data        ;
  output                                        mgr21__std__lane4_strm0_data_valid  ;

  input                                         std__mgr21__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane4_strm1_data        ;
  output                                        mgr21__std__lane4_strm1_data_valid  ;

  input                                         std__mgr21__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane5_strm0_data        ;
  output                                        mgr21__std__lane5_strm0_data_valid  ;

  input                                         std__mgr21__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane5_strm1_data        ;
  output                                        mgr21__std__lane5_strm1_data_valid  ;

  input                                         std__mgr21__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane6_strm0_data        ;
  output                                        mgr21__std__lane6_strm0_data_valid  ;

  input                                         std__mgr21__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane6_strm1_data        ;
  output                                        mgr21__std__lane6_strm1_data_valid  ;

  input                                         std__mgr21__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane7_strm0_data        ;
  output                                        mgr21__std__lane7_strm0_data_valid  ;

  input                                         std__mgr21__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane7_strm1_data        ;
  output                                        mgr21__std__lane7_strm1_data_valid  ;

  input                                         std__mgr21__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane8_strm0_data        ;
  output                                        mgr21__std__lane8_strm0_data_valid  ;

  input                                         std__mgr21__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane8_strm1_data        ;
  output                                        mgr21__std__lane8_strm1_data_valid  ;

  input                                         std__mgr21__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane9_strm0_data        ;
  output                                        mgr21__std__lane9_strm0_data_valid  ;

  input                                         std__mgr21__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane9_strm1_data        ;
  output                                        mgr21__std__lane9_strm1_data_valid  ;

  input                                         std__mgr21__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane10_strm0_data        ;
  output                                        mgr21__std__lane10_strm0_data_valid  ;

  input                                         std__mgr21__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane10_strm1_data        ;
  output                                        mgr21__std__lane10_strm1_data_valid  ;

  input                                         std__mgr21__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane11_strm0_data        ;
  output                                        mgr21__std__lane11_strm0_data_valid  ;

  input                                         std__mgr21__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane11_strm1_data        ;
  output                                        mgr21__std__lane11_strm1_data_valid  ;

  input                                         std__mgr21__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane12_strm0_data        ;
  output                                        mgr21__std__lane12_strm0_data_valid  ;

  input                                         std__mgr21__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane12_strm1_data        ;
  output                                        mgr21__std__lane12_strm1_data_valid  ;

  input                                         std__mgr21__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane13_strm0_data        ;
  output                                        mgr21__std__lane13_strm0_data_valid  ;

  input                                         std__mgr21__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane13_strm1_data        ;
  output                                        mgr21__std__lane13_strm1_data_valid  ;

  input                                         std__mgr21__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane14_strm0_data        ;
  output                                        mgr21__std__lane14_strm0_data_valid  ;

  input                                         std__mgr21__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane14_strm1_data        ;
  output                                        mgr21__std__lane14_strm1_data_valid  ;

  input                                         std__mgr21__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane15_strm0_data        ;
  output                                        mgr21__std__lane15_strm0_data_valid  ;

  input                                         std__mgr21__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane15_strm1_data        ;
  output                                        mgr21__std__lane15_strm1_data_valid  ;

  input                                         std__mgr21__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane16_strm0_data        ;
  output                                        mgr21__std__lane16_strm0_data_valid  ;

  input                                         std__mgr21__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane16_strm1_data        ;
  output                                        mgr21__std__lane16_strm1_data_valid  ;

  input                                         std__mgr21__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane17_strm0_data        ;
  output                                        mgr21__std__lane17_strm0_data_valid  ;

  input                                         std__mgr21__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane17_strm1_data        ;
  output                                        mgr21__std__lane17_strm1_data_valid  ;

  input                                         std__mgr21__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane18_strm0_data        ;
  output                                        mgr21__std__lane18_strm0_data_valid  ;

  input                                         std__mgr21__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane18_strm1_data        ;
  output                                        mgr21__std__lane18_strm1_data_valid  ;

  input                                         std__mgr21__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane19_strm0_data        ;
  output                                        mgr21__std__lane19_strm0_data_valid  ;

  input                                         std__mgr21__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane19_strm1_data        ;
  output                                        mgr21__std__lane19_strm1_data_valid  ;

  input                                         std__mgr21__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane20_strm0_data        ;
  output                                        mgr21__std__lane20_strm0_data_valid  ;

  input                                         std__mgr21__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane20_strm1_data        ;
  output                                        mgr21__std__lane20_strm1_data_valid  ;

  input                                         std__mgr21__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane21_strm0_data        ;
  output                                        mgr21__std__lane21_strm0_data_valid  ;

  input                                         std__mgr21__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane21_strm1_data        ;
  output                                        mgr21__std__lane21_strm1_data_valid  ;

  input                                         std__mgr21__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane22_strm0_data        ;
  output                                        mgr21__std__lane22_strm0_data_valid  ;

  input                                         std__mgr21__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane22_strm1_data        ;
  output                                        mgr21__std__lane22_strm1_data_valid  ;

  input                                         std__mgr21__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane23_strm0_data        ;
  output                                        mgr21__std__lane23_strm0_data_valid  ;

  input                                         std__mgr21__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane23_strm1_data        ;
  output                                        mgr21__std__lane23_strm1_data_valid  ;

  input                                         std__mgr21__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane24_strm0_data        ;
  output                                        mgr21__std__lane24_strm0_data_valid  ;

  input                                         std__mgr21__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane24_strm1_data        ;
  output                                        mgr21__std__lane24_strm1_data_valid  ;

  input                                         std__mgr21__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane25_strm0_data        ;
  output                                        mgr21__std__lane25_strm0_data_valid  ;

  input                                         std__mgr21__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane25_strm1_data        ;
  output                                        mgr21__std__lane25_strm1_data_valid  ;

  input                                         std__mgr21__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane26_strm0_data        ;
  output                                        mgr21__std__lane26_strm0_data_valid  ;

  input                                         std__mgr21__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane26_strm1_data        ;
  output                                        mgr21__std__lane26_strm1_data_valid  ;

  input                                         std__mgr21__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane27_strm0_data        ;
  output                                        mgr21__std__lane27_strm0_data_valid  ;

  input                                         std__mgr21__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane27_strm1_data        ;
  output                                        mgr21__std__lane27_strm1_data_valid  ;

  input                                         std__mgr21__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane28_strm0_data        ;
  output                                        mgr21__std__lane28_strm0_data_valid  ;

  input                                         std__mgr21__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane28_strm1_data        ;
  output                                        mgr21__std__lane28_strm1_data_valid  ;

  input                                         std__mgr21__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane29_strm0_data        ;
  output                                        mgr21__std__lane29_strm0_data_valid  ;

  input                                         std__mgr21__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane29_strm1_data        ;
  output                                        mgr21__std__lane29_strm1_data_valid  ;

  input                                         std__mgr21__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane30_strm0_data        ;
  output                                        mgr21__std__lane30_strm0_data_valid  ;

  input                                         std__mgr21__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane30_strm1_data        ;
  output                                        mgr21__std__lane30_strm1_data_valid  ;

  input                                         std__mgr21__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane31_strm0_data        ;
  output                                        mgr21__std__lane31_strm0_data_valid  ;

  input                                         std__mgr21__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane31_strm1_data        ;
  output                                        mgr21__std__lane31_strm1_data_valid  ;

  input                                         std__mgr22__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane0_strm0_data        ;
  output                                        mgr22__std__lane0_strm0_data_valid  ;

  input                                         std__mgr22__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane0_strm1_data        ;
  output                                        mgr22__std__lane0_strm1_data_valid  ;

  input                                         std__mgr22__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane1_strm0_data        ;
  output                                        mgr22__std__lane1_strm0_data_valid  ;

  input                                         std__mgr22__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane1_strm1_data        ;
  output                                        mgr22__std__lane1_strm1_data_valid  ;

  input                                         std__mgr22__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane2_strm0_data        ;
  output                                        mgr22__std__lane2_strm0_data_valid  ;

  input                                         std__mgr22__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane2_strm1_data        ;
  output                                        mgr22__std__lane2_strm1_data_valid  ;

  input                                         std__mgr22__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane3_strm0_data        ;
  output                                        mgr22__std__lane3_strm0_data_valid  ;

  input                                         std__mgr22__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane3_strm1_data        ;
  output                                        mgr22__std__lane3_strm1_data_valid  ;

  input                                         std__mgr22__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane4_strm0_data        ;
  output                                        mgr22__std__lane4_strm0_data_valid  ;

  input                                         std__mgr22__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane4_strm1_data        ;
  output                                        mgr22__std__lane4_strm1_data_valid  ;

  input                                         std__mgr22__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane5_strm0_data        ;
  output                                        mgr22__std__lane5_strm0_data_valid  ;

  input                                         std__mgr22__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane5_strm1_data        ;
  output                                        mgr22__std__lane5_strm1_data_valid  ;

  input                                         std__mgr22__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane6_strm0_data        ;
  output                                        mgr22__std__lane6_strm0_data_valid  ;

  input                                         std__mgr22__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane6_strm1_data        ;
  output                                        mgr22__std__lane6_strm1_data_valid  ;

  input                                         std__mgr22__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane7_strm0_data        ;
  output                                        mgr22__std__lane7_strm0_data_valid  ;

  input                                         std__mgr22__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane7_strm1_data        ;
  output                                        mgr22__std__lane7_strm1_data_valid  ;

  input                                         std__mgr22__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane8_strm0_data        ;
  output                                        mgr22__std__lane8_strm0_data_valid  ;

  input                                         std__mgr22__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane8_strm1_data        ;
  output                                        mgr22__std__lane8_strm1_data_valid  ;

  input                                         std__mgr22__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane9_strm0_data        ;
  output                                        mgr22__std__lane9_strm0_data_valid  ;

  input                                         std__mgr22__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane9_strm1_data        ;
  output                                        mgr22__std__lane9_strm1_data_valid  ;

  input                                         std__mgr22__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane10_strm0_data        ;
  output                                        mgr22__std__lane10_strm0_data_valid  ;

  input                                         std__mgr22__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane10_strm1_data        ;
  output                                        mgr22__std__lane10_strm1_data_valid  ;

  input                                         std__mgr22__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane11_strm0_data        ;
  output                                        mgr22__std__lane11_strm0_data_valid  ;

  input                                         std__mgr22__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane11_strm1_data        ;
  output                                        mgr22__std__lane11_strm1_data_valid  ;

  input                                         std__mgr22__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane12_strm0_data        ;
  output                                        mgr22__std__lane12_strm0_data_valid  ;

  input                                         std__mgr22__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane12_strm1_data        ;
  output                                        mgr22__std__lane12_strm1_data_valid  ;

  input                                         std__mgr22__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane13_strm0_data        ;
  output                                        mgr22__std__lane13_strm0_data_valid  ;

  input                                         std__mgr22__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane13_strm1_data        ;
  output                                        mgr22__std__lane13_strm1_data_valid  ;

  input                                         std__mgr22__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane14_strm0_data        ;
  output                                        mgr22__std__lane14_strm0_data_valid  ;

  input                                         std__mgr22__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane14_strm1_data        ;
  output                                        mgr22__std__lane14_strm1_data_valid  ;

  input                                         std__mgr22__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane15_strm0_data        ;
  output                                        mgr22__std__lane15_strm0_data_valid  ;

  input                                         std__mgr22__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane15_strm1_data        ;
  output                                        mgr22__std__lane15_strm1_data_valid  ;

  input                                         std__mgr22__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane16_strm0_data        ;
  output                                        mgr22__std__lane16_strm0_data_valid  ;

  input                                         std__mgr22__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane16_strm1_data        ;
  output                                        mgr22__std__lane16_strm1_data_valid  ;

  input                                         std__mgr22__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane17_strm0_data        ;
  output                                        mgr22__std__lane17_strm0_data_valid  ;

  input                                         std__mgr22__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane17_strm1_data        ;
  output                                        mgr22__std__lane17_strm1_data_valid  ;

  input                                         std__mgr22__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane18_strm0_data        ;
  output                                        mgr22__std__lane18_strm0_data_valid  ;

  input                                         std__mgr22__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane18_strm1_data        ;
  output                                        mgr22__std__lane18_strm1_data_valid  ;

  input                                         std__mgr22__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane19_strm0_data        ;
  output                                        mgr22__std__lane19_strm0_data_valid  ;

  input                                         std__mgr22__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane19_strm1_data        ;
  output                                        mgr22__std__lane19_strm1_data_valid  ;

  input                                         std__mgr22__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane20_strm0_data        ;
  output                                        mgr22__std__lane20_strm0_data_valid  ;

  input                                         std__mgr22__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane20_strm1_data        ;
  output                                        mgr22__std__lane20_strm1_data_valid  ;

  input                                         std__mgr22__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane21_strm0_data        ;
  output                                        mgr22__std__lane21_strm0_data_valid  ;

  input                                         std__mgr22__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane21_strm1_data        ;
  output                                        mgr22__std__lane21_strm1_data_valid  ;

  input                                         std__mgr22__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane22_strm0_data        ;
  output                                        mgr22__std__lane22_strm0_data_valid  ;

  input                                         std__mgr22__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane22_strm1_data        ;
  output                                        mgr22__std__lane22_strm1_data_valid  ;

  input                                         std__mgr22__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane23_strm0_data        ;
  output                                        mgr22__std__lane23_strm0_data_valid  ;

  input                                         std__mgr22__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane23_strm1_data        ;
  output                                        mgr22__std__lane23_strm1_data_valid  ;

  input                                         std__mgr22__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane24_strm0_data        ;
  output                                        mgr22__std__lane24_strm0_data_valid  ;

  input                                         std__mgr22__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane24_strm1_data        ;
  output                                        mgr22__std__lane24_strm1_data_valid  ;

  input                                         std__mgr22__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane25_strm0_data        ;
  output                                        mgr22__std__lane25_strm0_data_valid  ;

  input                                         std__mgr22__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane25_strm1_data        ;
  output                                        mgr22__std__lane25_strm1_data_valid  ;

  input                                         std__mgr22__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane26_strm0_data        ;
  output                                        mgr22__std__lane26_strm0_data_valid  ;

  input                                         std__mgr22__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane26_strm1_data        ;
  output                                        mgr22__std__lane26_strm1_data_valid  ;

  input                                         std__mgr22__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane27_strm0_data        ;
  output                                        mgr22__std__lane27_strm0_data_valid  ;

  input                                         std__mgr22__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane27_strm1_data        ;
  output                                        mgr22__std__lane27_strm1_data_valid  ;

  input                                         std__mgr22__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane28_strm0_data        ;
  output                                        mgr22__std__lane28_strm0_data_valid  ;

  input                                         std__mgr22__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane28_strm1_data        ;
  output                                        mgr22__std__lane28_strm1_data_valid  ;

  input                                         std__mgr22__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane29_strm0_data        ;
  output                                        mgr22__std__lane29_strm0_data_valid  ;

  input                                         std__mgr22__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane29_strm1_data        ;
  output                                        mgr22__std__lane29_strm1_data_valid  ;

  input                                         std__mgr22__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane30_strm0_data        ;
  output                                        mgr22__std__lane30_strm0_data_valid  ;

  input                                         std__mgr22__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane30_strm1_data        ;
  output                                        mgr22__std__lane30_strm1_data_valid  ;

  input                                         std__mgr22__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane31_strm0_data        ;
  output                                        mgr22__std__lane31_strm0_data_valid  ;

  input                                         std__mgr22__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane31_strm1_data        ;
  output                                        mgr22__std__lane31_strm1_data_valid  ;

  input                                         std__mgr23__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane0_strm0_data        ;
  output                                        mgr23__std__lane0_strm0_data_valid  ;

  input                                         std__mgr23__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane0_strm1_data        ;
  output                                        mgr23__std__lane0_strm1_data_valid  ;

  input                                         std__mgr23__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane1_strm0_data        ;
  output                                        mgr23__std__lane1_strm0_data_valid  ;

  input                                         std__mgr23__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane1_strm1_data        ;
  output                                        mgr23__std__lane1_strm1_data_valid  ;

  input                                         std__mgr23__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane2_strm0_data        ;
  output                                        mgr23__std__lane2_strm0_data_valid  ;

  input                                         std__mgr23__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane2_strm1_data        ;
  output                                        mgr23__std__lane2_strm1_data_valid  ;

  input                                         std__mgr23__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane3_strm0_data        ;
  output                                        mgr23__std__lane3_strm0_data_valid  ;

  input                                         std__mgr23__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane3_strm1_data        ;
  output                                        mgr23__std__lane3_strm1_data_valid  ;

  input                                         std__mgr23__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane4_strm0_data        ;
  output                                        mgr23__std__lane4_strm0_data_valid  ;

  input                                         std__mgr23__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane4_strm1_data        ;
  output                                        mgr23__std__lane4_strm1_data_valid  ;

  input                                         std__mgr23__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane5_strm0_data        ;
  output                                        mgr23__std__lane5_strm0_data_valid  ;

  input                                         std__mgr23__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane5_strm1_data        ;
  output                                        mgr23__std__lane5_strm1_data_valid  ;

  input                                         std__mgr23__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane6_strm0_data        ;
  output                                        mgr23__std__lane6_strm0_data_valid  ;

  input                                         std__mgr23__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane6_strm1_data        ;
  output                                        mgr23__std__lane6_strm1_data_valid  ;

  input                                         std__mgr23__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane7_strm0_data        ;
  output                                        mgr23__std__lane7_strm0_data_valid  ;

  input                                         std__mgr23__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane7_strm1_data        ;
  output                                        mgr23__std__lane7_strm1_data_valid  ;

  input                                         std__mgr23__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane8_strm0_data        ;
  output                                        mgr23__std__lane8_strm0_data_valid  ;

  input                                         std__mgr23__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane8_strm1_data        ;
  output                                        mgr23__std__lane8_strm1_data_valid  ;

  input                                         std__mgr23__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane9_strm0_data        ;
  output                                        mgr23__std__lane9_strm0_data_valid  ;

  input                                         std__mgr23__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane9_strm1_data        ;
  output                                        mgr23__std__lane9_strm1_data_valid  ;

  input                                         std__mgr23__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane10_strm0_data        ;
  output                                        mgr23__std__lane10_strm0_data_valid  ;

  input                                         std__mgr23__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane10_strm1_data        ;
  output                                        mgr23__std__lane10_strm1_data_valid  ;

  input                                         std__mgr23__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane11_strm0_data        ;
  output                                        mgr23__std__lane11_strm0_data_valid  ;

  input                                         std__mgr23__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane11_strm1_data        ;
  output                                        mgr23__std__lane11_strm1_data_valid  ;

  input                                         std__mgr23__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane12_strm0_data        ;
  output                                        mgr23__std__lane12_strm0_data_valid  ;

  input                                         std__mgr23__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane12_strm1_data        ;
  output                                        mgr23__std__lane12_strm1_data_valid  ;

  input                                         std__mgr23__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane13_strm0_data        ;
  output                                        mgr23__std__lane13_strm0_data_valid  ;

  input                                         std__mgr23__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane13_strm1_data        ;
  output                                        mgr23__std__lane13_strm1_data_valid  ;

  input                                         std__mgr23__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane14_strm0_data        ;
  output                                        mgr23__std__lane14_strm0_data_valid  ;

  input                                         std__mgr23__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane14_strm1_data        ;
  output                                        mgr23__std__lane14_strm1_data_valid  ;

  input                                         std__mgr23__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane15_strm0_data        ;
  output                                        mgr23__std__lane15_strm0_data_valid  ;

  input                                         std__mgr23__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane15_strm1_data        ;
  output                                        mgr23__std__lane15_strm1_data_valid  ;

  input                                         std__mgr23__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane16_strm0_data        ;
  output                                        mgr23__std__lane16_strm0_data_valid  ;

  input                                         std__mgr23__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane16_strm1_data        ;
  output                                        mgr23__std__lane16_strm1_data_valid  ;

  input                                         std__mgr23__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane17_strm0_data        ;
  output                                        mgr23__std__lane17_strm0_data_valid  ;

  input                                         std__mgr23__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane17_strm1_data        ;
  output                                        mgr23__std__lane17_strm1_data_valid  ;

  input                                         std__mgr23__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane18_strm0_data        ;
  output                                        mgr23__std__lane18_strm0_data_valid  ;

  input                                         std__mgr23__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane18_strm1_data        ;
  output                                        mgr23__std__lane18_strm1_data_valid  ;

  input                                         std__mgr23__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane19_strm0_data        ;
  output                                        mgr23__std__lane19_strm0_data_valid  ;

  input                                         std__mgr23__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane19_strm1_data        ;
  output                                        mgr23__std__lane19_strm1_data_valid  ;

  input                                         std__mgr23__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane20_strm0_data        ;
  output                                        mgr23__std__lane20_strm0_data_valid  ;

  input                                         std__mgr23__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane20_strm1_data        ;
  output                                        mgr23__std__lane20_strm1_data_valid  ;

  input                                         std__mgr23__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane21_strm0_data        ;
  output                                        mgr23__std__lane21_strm0_data_valid  ;

  input                                         std__mgr23__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane21_strm1_data        ;
  output                                        mgr23__std__lane21_strm1_data_valid  ;

  input                                         std__mgr23__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane22_strm0_data        ;
  output                                        mgr23__std__lane22_strm0_data_valid  ;

  input                                         std__mgr23__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane22_strm1_data        ;
  output                                        mgr23__std__lane22_strm1_data_valid  ;

  input                                         std__mgr23__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane23_strm0_data        ;
  output                                        mgr23__std__lane23_strm0_data_valid  ;

  input                                         std__mgr23__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane23_strm1_data        ;
  output                                        mgr23__std__lane23_strm1_data_valid  ;

  input                                         std__mgr23__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane24_strm0_data        ;
  output                                        mgr23__std__lane24_strm0_data_valid  ;

  input                                         std__mgr23__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane24_strm1_data        ;
  output                                        mgr23__std__lane24_strm1_data_valid  ;

  input                                         std__mgr23__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane25_strm0_data        ;
  output                                        mgr23__std__lane25_strm0_data_valid  ;

  input                                         std__mgr23__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane25_strm1_data        ;
  output                                        mgr23__std__lane25_strm1_data_valid  ;

  input                                         std__mgr23__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane26_strm0_data        ;
  output                                        mgr23__std__lane26_strm0_data_valid  ;

  input                                         std__mgr23__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane26_strm1_data        ;
  output                                        mgr23__std__lane26_strm1_data_valid  ;

  input                                         std__mgr23__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane27_strm0_data        ;
  output                                        mgr23__std__lane27_strm0_data_valid  ;

  input                                         std__mgr23__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane27_strm1_data        ;
  output                                        mgr23__std__lane27_strm1_data_valid  ;

  input                                         std__mgr23__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane28_strm0_data        ;
  output                                        mgr23__std__lane28_strm0_data_valid  ;

  input                                         std__mgr23__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane28_strm1_data        ;
  output                                        mgr23__std__lane28_strm1_data_valid  ;

  input                                         std__mgr23__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane29_strm0_data        ;
  output                                        mgr23__std__lane29_strm0_data_valid  ;

  input                                         std__mgr23__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane29_strm1_data        ;
  output                                        mgr23__std__lane29_strm1_data_valid  ;

  input                                         std__mgr23__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane30_strm0_data        ;
  output                                        mgr23__std__lane30_strm0_data_valid  ;

  input                                         std__mgr23__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane30_strm1_data        ;
  output                                        mgr23__std__lane30_strm1_data_valid  ;

  input                                         std__mgr23__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane31_strm0_data        ;
  output                                        mgr23__std__lane31_strm0_data_valid  ;

  input                                         std__mgr23__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane31_strm1_data        ;
  output                                        mgr23__std__lane31_strm1_data_valid  ;

  input                                         std__mgr24__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane0_strm0_data        ;
  output                                        mgr24__std__lane0_strm0_data_valid  ;

  input                                         std__mgr24__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane0_strm1_data        ;
  output                                        mgr24__std__lane0_strm1_data_valid  ;

  input                                         std__mgr24__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane1_strm0_data        ;
  output                                        mgr24__std__lane1_strm0_data_valid  ;

  input                                         std__mgr24__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane1_strm1_data        ;
  output                                        mgr24__std__lane1_strm1_data_valid  ;

  input                                         std__mgr24__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane2_strm0_data        ;
  output                                        mgr24__std__lane2_strm0_data_valid  ;

  input                                         std__mgr24__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane2_strm1_data        ;
  output                                        mgr24__std__lane2_strm1_data_valid  ;

  input                                         std__mgr24__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane3_strm0_data        ;
  output                                        mgr24__std__lane3_strm0_data_valid  ;

  input                                         std__mgr24__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane3_strm1_data        ;
  output                                        mgr24__std__lane3_strm1_data_valid  ;

  input                                         std__mgr24__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane4_strm0_data        ;
  output                                        mgr24__std__lane4_strm0_data_valid  ;

  input                                         std__mgr24__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane4_strm1_data        ;
  output                                        mgr24__std__lane4_strm1_data_valid  ;

  input                                         std__mgr24__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane5_strm0_data        ;
  output                                        mgr24__std__lane5_strm0_data_valid  ;

  input                                         std__mgr24__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane5_strm1_data        ;
  output                                        mgr24__std__lane5_strm1_data_valid  ;

  input                                         std__mgr24__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane6_strm0_data        ;
  output                                        mgr24__std__lane6_strm0_data_valid  ;

  input                                         std__mgr24__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane6_strm1_data        ;
  output                                        mgr24__std__lane6_strm1_data_valid  ;

  input                                         std__mgr24__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane7_strm0_data        ;
  output                                        mgr24__std__lane7_strm0_data_valid  ;

  input                                         std__mgr24__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane7_strm1_data        ;
  output                                        mgr24__std__lane7_strm1_data_valid  ;

  input                                         std__mgr24__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane8_strm0_data        ;
  output                                        mgr24__std__lane8_strm0_data_valid  ;

  input                                         std__mgr24__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane8_strm1_data        ;
  output                                        mgr24__std__lane8_strm1_data_valid  ;

  input                                         std__mgr24__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane9_strm0_data        ;
  output                                        mgr24__std__lane9_strm0_data_valid  ;

  input                                         std__mgr24__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane9_strm1_data        ;
  output                                        mgr24__std__lane9_strm1_data_valid  ;

  input                                         std__mgr24__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane10_strm0_data        ;
  output                                        mgr24__std__lane10_strm0_data_valid  ;

  input                                         std__mgr24__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane10_strm1_data        ;
  output                                        mgr24__std__lane10_strm1_data_valid  ;

  input                                         std__mgr24__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane11_strm0_data        ;
  output                                        mgr24__std__lane11_strm0_data_valid  ;

  input                                         std__mgr24__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane11_strm1_data        ;
  output                                        mgr24__std__lane11_strm1_data_valid  ;

  input                                         std__mgr24__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane12_strm0_data        ;
  output                                        mgr24__std__lane12_strm0_data_valid  ;

  input                                         std__mgr24__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane12_strm1_data        ;
  output                                        mgr24__std__lane12_strm1_data_valid  ;

  input                                         std__mgr24__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane13_strm0_data        ;
  output                                        mgr24__std__lane13_strm0_data_valid  ;

  input                                         std__mgr24__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane13_strm1_data        ;
  output                                        mgr24__std__lane13_strm1_data_valid  ;

  input                                         std__mgr24__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane14_strm0_data        ;
  output                                        mgr24__std__lane14_strm0_data_valid  ;

  input                                         std__mgr24__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane14_strm1_data        ;
  output                                        mgr24__std__lane14_strm1_data_valid  ;

  input                                         std__mgr24__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane15_strm0_data        ;
  output                                        mgr24__std__lane15_strm0_data_valid  ;

  input                                         std__mgr24__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane15_strm1_data        ;
  output                                        mgr24__std__lane15_strm1_data_valid  ;

  input                                         std__mgr24__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane16_strm0_data        ;
  output                                        mgr24__std__lane16_strm0_data_valid  ;

  input                                         std__mgr24__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane16_strm1_data        ;
  output                                        mgr24__std__lane16_strm1_data_valid  ;

  input                                         std__mgr24__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane17_strm0_data        ;
  output                                        mgr24__std__lane17_strm0_data_valid  ;

  input                                         std__mgr24__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane17_strm1_data        ;
  output                                        mgr24__std__lane17_strm1_data_valid  ;

  input                                         std__mgr24__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane18_strm0_data        ;
  output                                        mgr24__std__lane18_strm0_data_valid  ;

  input                                         std__mgr24__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane18_strm1_data        ;
  output                                        mgr24__std__lane18_strm1_data_valid  ;

  input                                         std__mgr24__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane19_strm0_data        ;
  output                                        mgr24__std__lane19_strm0_data_valid  ;

  input                                         std__mgr24__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane19_strm1_data        ;
  output                                        mgr24__std__lane19_strm1_data_valid  ;

  input                                         std__mgr24__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane20_strm0_data        ;
  output                                        mgr24__std__lane20_strm0_data_valid  ;

  input                                         std__mgr24__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane20_strm1_data        ;
  output                                        mgr24__std__lane20_strm1_data_valid  ;

  input                                         std__mgr24__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane21_strm0_data        ;
  output                                        mgr24__std__lane21_strm0_data_valid  ;

  input                                         std__mgr24__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane21_strm1_data        ;
  output                                        mgr24__std__lane21_strm1_data_valid  ;

  input                                         std__mgr24__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane22_strm0_data        ;
  output                                        mgr24__std__lane22_strm0_data_valid  ;

  input                                         std__mgr24__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane22_strm1_data        ;
  output                                        mgr24__std__lane22_strm1_data_valid  ;

  input                                         std__mgr24__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane23_strm0_data        ;
  output                                        mgr24__std__lane23_strm0_data_valid  ;

  input                                         std__mgr24__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane23_strm1_data        ;
  output                                        mgr24__std__lane23_strm1_data_valid  ;

  input                                         std__mgr24__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane24_strm0_data        ;
  output                                        mgr24__std__lane24_strm0_data_valid  ;

  input                                         std__mgr24__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane24_strm1_data        ;
  output                                        mgr24__std__lane24_strm1_data_valid  ;

  input                                         std__mgr24__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane25_strm0_data        ;
  output                                        mgr24__std__lane25_strm0_data_valid  ;

  input                                         std__mgr24__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane25_strm1_data        ;
  output                                        mgr24__std__lane25_strm1_data_valid  ;

  input                                         std__mgr24__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane26_strm0_data        ;
  output                                        mgr24__std__lane26_strm0_data_valid  ;

  input                                         std__mgr24__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane26_strm1_data        ;
  output                                        mgr24__std__lane26_strm1_data_valid  ;

  input                                         std__mgr24__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane27_strm0_data        ;
  output                                        mgr24__std__lane27_strm0_data_valid  ;

  input                                         std__mgr24__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane27_strm1_data        ;
  output                                        mgr24__std__lane27_strm1_data_valid  ;

  input                                         std__mgr24__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane28_strm0_data        ;
  output                                        mgr24__std__lane28_strm0_data_valid  ;

  input                                         std__mgr24__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane28_strm1_data        ;
  output                                        mgr24__std__lane28_strm1_data_valid  ;

  input                                         std__mgr24__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane29_strm0_data        ;
  output                                        mgr24__std__lane29_strm0_data_valid  ;

  input                                         std__mgr24__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane29_strm1_data        ;
  output                                        mgr24__std__lane29_strm1_data_valid  ;

  input                                         std__mgr24__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane30_strm0_data        ;
  output                                        mgr24__std__lane30_strm0_data_valid  ;

  input                                         std__mgr24__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane30_strm1_data        ;
  output                                        mgr24__std__lane30_strm1_data_valid  ;

  input                                         std__mgr24__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane31_strm0_data        ;
  output                                        mgr24__std__lane31_strm0_data_valid  ;

  input                                         std__mgr24__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane31_strm1_data        ;
  output                                        mgr24__std__lane31_strm1_data_valid  ;

  input                                         std__mgr25__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane0_strm0_data        ;
  output                                        mgr25__std__lane0_strm0_data_valid  ;

  input                                         std__mgr25__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane0_strm1_data        ;
  output                                        mgr25__std__lane0_strm1_data_valid  ;

  input                                         std__mgr25__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane1_strm0_data        ;
  output                                        mgr25__std__lane1_strm0_data_valid  ;

  input                                         std__mgr25__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane1_strm1_data        ;
  output                                        mgr25__std__lane1_strm1_data_valid  ;

  input                                         std__mgr25__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane2_strm0_data        ;
  output                                        mgr25__std__lane2_strm0_data_valid  ;

  input                                         std__mgr25__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane2_strm1_data        ;
  output                                        mgr25__std__lane2_strm1_data_valid  ;

  input                                         std__mgr25__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane3_strm0_data        ;
  output                                        mgr25__std__lane3_strm0_data_valid  ;

  input                                         std__mgr25__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane3_strm1_data        ;
  output                                        mgr25__std__lane3_strm1_data_valid  ;

  input                                         std__mgr25__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane4_strm0_data        ;
  output                                        mgr25__std__lane4_strm0_data_valid  ;

  input                                         std__mgr25__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane4_strm1_data        ;
  output                                        mgr25__std__lane4_strm1_data_valid  ;

  input                                         std__mgr25__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane5_strm0_data        ;
  output                                        mgr25__std__lane5_strm0_data_valid  ;

  input                                         std__mgr25__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane5_strm1_data        ;
  output                                        mgr25__std__lane5_strm1_data_valid  ;

  input                                         std__mgr25__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane6_strm0_data        ;
  output                                        mgr25__std__lane6_strm0_data_valid  ;

  input                                         std__mgr25__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane6_strm1_data        ;
  output                                        mgr25__std__lane6_strm1_data_valid  ;

  input                                         std__mgr25__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane7_strm0_data        ;
  output                                        mgr25__std__lane7_strm0_data_valid  ;

  input                                         std__mgr25__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane7_strm1_data        ;
  output                                        mgr25__std__lane7_strm1_data_valid  ;

  input                                         std__mgr25__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane8_strm0_data        ;
  output                                        mgr25__std__lane8_strm0_data_valid  ;

  input                                         std__mgr25__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane8_strm1_data        ;
  output                                        mgr25__std__lane8_strm1_data_valid  ;

  input                                         std__mgr25__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane9_strm0_data        ;
  output                                        mgr25__std__lane9_strm0_data_valid  ;

  input                                         std__mgr25__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane9_strm1_data        ;
  output                                        mgr25__std__lane9_strm1_data_valid  ;

  input                                         std__mgr25__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane10_strm0_data        ;
  output                                        mgr25__std__lane10_strm0_data_valid  ;

  input                                         std__mgr25__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane10_strm1_data        ;
  output                                        mgr25__std__lane10_strm1_data_valid  ;

  input                                         std__mgr25__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane11_strm0_data        ;
  output                                        mgr25__std__lane11_strm0_data_valid  ;

  input                                         std__mgr25__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane11_strm1_data        ;
  output                                        mgr25__std__lane11_strm1_data_valid  ;

  input                                         std__mgr25__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane12_strm0_data        ;
  output                                        mgr25__std__lane12_strm0_data_valid  ;

  input                                         std__mgr25__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane12_strm1_data        ;
  output                                        mgr25__std__lane12_strm1_data_valid  ;

  input                                         std__mgr25__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane13_strm0_data        ;
  output                                        mgr25__std__lane13_strm0_data_valid  ;

  input                                         std__mgr25__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane13_strm1_data        ;
  output                                        mgr25__std__lane13_strm1_data_valid  ;

  input                                         std__mgr25__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane14_strm0_data        ;
  output                                        mgr25__std__lane14_strm0_data_valid  ;

  input                                         std__mgr25__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane14_strm1_data        ;
  output                                        mgr25__std__lane14_strm1_data_valid  ;

  input                                         std__mgr25__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane15_strm0_data        ;
  output                                        mgr25__std__lane15_strm0_data_valid  ;

  input                                         std__mgr25__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane15_strm1_data        ;
  output                                        mgr25__std__lane15_strm1_data_valid  ;

  input                                         std__mgr25__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane16_strm0_data        ;
  output                                        mgr25__std__lane16_strm0_data_valid  ;

  input                                         std__mgr25__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane16_strm1_data        ;
  output                                        mgr25__std__lane16_strm1_data_valid  ;

  input                                         std__mgr25__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane17_strm0_data        ;
  output                                        mgr25__std__lane17_strm0_data_valid  ;

  input                                         std__mgr25__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane17_strm1_data        ;
  output                                        mgr25__std__lane17_strm1_data_valid  ;

  input                                         std__mgr25__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane18_strm0_data        ;
  output                                        mgr25__std__lane18_strm0_data_valid  ;

  input                                         std__mgr25__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane18_strm1_data        ;
  output                                        mgr25__std__lane18_strm1_data_valid  ;

  input                                         std__mgr25__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane19_strm0_data        ;
  output                                        mgr25__std__lane19_strm0_data_valid  ;

  input                                         std__mgr25__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane19_strm1_data        ;
  output                                        mgr25__std__lane19_strm1_data_valid  ;

  input                                         std__mgr25__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane20_strm0_data        ;
  output                                        mgr25__std__lane20_strm0_data_valid  ;

  input                                         std__mgr25__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane20_strm1_data        ;
  output                                        mgr25__std__lane20_strm1_data_valid  ;

  input                                         std__mgr25__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane21_strm0_data        ;
  output                                        mgr25__std__lane21_strm0_data_valid  ;

  input                                         std__mgr25__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane21_strm1_data        ;
  output                                        mgr25__std__lane21_strm1_data_valid  ;

  input                                         std__mgr25__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane22_strm0_data        ;
  output                                        mgr25__std__lane22_strm0_data_valid  ;

  input                                         std__mgr25__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane22_strm1_data        ;
  output                                        mgr25__std__lane22_strm1_data_valid  ;

  input                                         std__mgr25__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane23_strm0_data        ;
  output                                        mgr25__std__lane23_strm0_data_valid  ;

  input                                         std__mgr25__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane23_strm1_data        ;
  output                                        mgr25__std__lane23_strm1_data_valid  ;

  input                                         std__mgr25__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane24_strm0_data        ;
  output                                        mgr25__std__lane24_strm0_data_valid  ;

  input                                         std__mgr25__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane24_strm1_data        ;
  output                                        mgr25__std__lane24_strm1_data_valid  ;

  input                                         std__mgr25__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane25_strm0_data        ;
  output                                        mgr25__std__lane25_strm0_data_valid  ;

  input                                         std__mgr25__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane25_strm1_data        ;
  output                                        mgr25__std__lane25_strm1_data_valid  ;

  input                                         std__mgr25__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane26_strm0_data        ;
  output                                        mgr25__std__lane26_strm0_data_valid  ;

  input                                         std__mgr25__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane26_strm1_data        ;
  output                                        mgr25__std__lane26_strm1_data_valid  ;

  input                                         std__mgr25__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane27_strm0_data        ;
  output                                        mgr25__std__lane27_strm0_data_valid  ;

  input                                         std__mgr25__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane27_strm1_data        ;
  output                                        mgr25__std__lane27_strm1_data_valid  ;

  input                                         std__mgr25__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane28_strm0_data        ;
  output                                        mgr25__std__lane28_strm0_data_valid  ;

  input                                         std__mgr25__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane28_strm1_data        ;
  output                                        mgr25__std__lane28_strm1_data_valid  ;

  input                                         std__mgr25__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane29_strm0_data        ;
  output                                        mgr25__std__lane29_strm0_data_valid  ;

  input                                         std__mgr25__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane29_strm1_data        ;
  output                                        mgr25__std__lane29_strm1_data_valid  ;

  input                                         std__mgr25__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane30_strm0_data        ;
  output                                        mgr25__std__lane30_strm0_data_valid  ;

  input                                         std__mgr25__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane30_strm1_data        ;
  output                                        mgr25__std__lane30_strm1_data_valid  ;

  input                                         std__mgr25__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane31_strm0_data        ;
  output                                        mgr25__std__lane31_strm0_data_valid  ;

  input                                         std__mgr25__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane31_strm1_data        ;
  output                                        mgr25__std__lane31_strm1_data_valid  ;

  input                                         std__mgr26__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane0_strm0_data        ;
  output                                        mgr26__std__lane0_strm0_data_valid  ;

  input                                         std__mgr26__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane0_strm1_data        ;
  output                                        mgr26__std__lane0_strm1_data_valid  ;

  input                                         std__mgr26__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane1_strm0_data        ;
  output                                        mgr26__std__lane1_strm0_data_valid  ;

  input                                         std__mgr26__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane1_strm1_data        ;
  output                                        mgr26__std__lane1_strm1_data_valid  ;

  input                                         std__mgr26__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane2_strm0_data        ;
  output                                        mgr26__std__lane2_strm0_data_valid  ;

  input                                         std__mgr26__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane2_strm1_data        ;
  output                                        mgr26__std__lane2_strm1_data_valid  ;

  input                                         std__mgr26__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane3_strm0_data        ;
  output                                        mgr26__std__lane3_strm0_data_valid  ;

  input                                         std__mgr26__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane3_strm1_data        ;
  output                                        mgr26__std__lane3_strm1_data_valid  ;

  input                                         std__mgr26__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane4_strm0_data        ;
  output                                        mgr26__std__lane4_strm0_data_valid  ;

  input                                         std__mgr26__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane4_strm1_data        ;
  output                                        mgr26__std__lane4_strm1_data_valid  ;

  input                                         std__mgr26__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane5_strm0_data        ;
  output                                        mgr26__std__lane5_strm0_data_valid  ;

  input                                         std__mgr26__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane5_strm1_data        ;
  output                                        mgr26__std__lane5_strm1_data_valid  ;

  input                                         std__mgr26__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane6_strm0_data        ;
  output                                        mgr26__std__lane6_strm0_data_valid  ;

  input                                         std__mgr26__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane6_strm1_data        ;
  output                                        mgr26__std__lane6_strm1_data_valid  ;

  input                                         std__mgr26__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane7_strm0_data        ;
  output                                        mgr26__std__lane7_strm0_data_valid  ;

  input                                         std__mgr26__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane7_strm1_data        ;
  output                                        mgr26__std__lane7_strm1_data_valid  ;

  input                                         std__mgr26__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane8_strm0_data        ;
  output                                        mgr26__std__lane8_strm0_data_valid  ;

  input                                         std__mgr26__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane8_strm1_data        ;
  output                                        mgr26__std__lane8_strm1_data_valid  ;

  input                                         std__mgr26__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane9_strm0_data        ;
  output                                        mgr26__std__lane9_strm0_data_valid  ;

  input                                         std__mgr26__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane9_strm1_data        ;
  output                                        mgr26__std__lane9_strm1_data_valid  ;

  input                                         std__mgr26__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane10_strm0_data        ;
  output                                        mgr26__std__lane10_strm0_data_valid  ;

  input                                         std__mgr26__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane10_strm1_data        ;
  output                                        mgr26__std__lane10_strm1_data_valid  ;

  input                                         std__mgr26__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane11_strm0_data        ;
  output                                        mgr26__std__lane11_strm0_data_valid  ;

  input                                         std__mgr26__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane11_strm1_data        ;
  output                                        mgr26__std__lane11_strm1_data_valid  ;

  input                                         std__mgr26__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane12_strm0_data        ;
  output                                        mgr26__std__lane12_strm0_data_valid  ;

  input                                         std__mgr26__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane12_strm1_data        ;
  output                                        mgr26__std__lane12_strm1_data_valid  ;

  input                                         std__mgr26__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane13_strm0_data        ;
  output                                        mgr26__std__lane13_strm0_data_valid  ;

  input                                         std__mgr26__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane13_strm1_data        ;
  output                                        mgr26__std__lane13_strm1_data_valid  ;

  input                                         std__mgr26__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane14_strm0_data        ;
  output                                        mgr26__std__lane14_strm0_data_valid  ;

  input                                         std__mgr26__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane14_strm1_data        ;
  output                                        mgr26__std__lane14_strm1_data_valid  ;

  input                                         std__mgr26__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane15_strm0_data        ;
  output                                        mgr26__std__lane15_strm0_data_valid  ;

  input                                         std__mgr26__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane15_strm1_data        ;
  output                                        mgr26__std__lane15_strm1_data_valid  ;

  input                                         std__mgr26__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane16_strm0_data        ;
  output                                        mgr26__std__lane16_strm0_data_valid  ;

  input                                         std__mgr26__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane16_strm1_data        ;
  output                                        mgr26__std__lane16_strm1_data_valid  ;

  input                                         std__mgr26__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane17_strm0_data        ;
  output                                        mgr26__std__lane17_strm0_data_valid  ;

  input                                         std__mgr26__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane17_strm1_data        ;
  output                                        mgr26__std__lane17_strm1_data_valid  ;

  input                                         std__mgr26__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane18_strm0_data        ;
  output                                        mgr26__std__lane18_strm0_data_valid  ;

  input                                         std__mgr26__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane18_strm1_data        ;
  output                                        mgr26__std__lane18_strm1_data_valid  ;

  input                                         std__mgr26__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane19_strm0_data        ;
  output                                        mgr26__std__lane19_strm0_data_valid  ;

  input                                         std__mgr26__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane19_strm1_data        ;
  output                                        mgr26__std__lane19_strm1_data_valid  ;

  input                                         std__mgr26__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane20_strm0_data        ;
  output                                        mgr26__std__lane20_strm0_data_valid  ;

  input                                         std__mgr26__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane20_strm1_data        ;
  output                                        mgr26__std__lane20_strm1_data_valid  ;

  input                                         std__mgr26__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane21_strm0_data        ;
  output                                        mgr26__std__lane21_strm0_data_valid  ;

  input                                         std__mgr26__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane21_strm1_data        ;
  output                                        mgr26__std__lane21_strm1_data_valid  ;

  input                                         std__mgr26__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane22_strm0_data        ;
  output                                        mgr26__std__lane22_strm0_data_valid  ;

  input                                         std__mgr26__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane22_strm1_data        ;
  output                                        mgr26__std__lane22_strm1_data_valid  ;

  input                                         std__mgr26__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane23_strm0_data        ;
  output                                        mgr26__std__lane23_strm0_data_valid  ;

  input                                         std__mgr26__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane23_strm1_data        ;
  output                                        mgr26__std__lane23_strm1_data_valid  ;

  input                                         std__mgr26__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane24_strm0_data        ;
  output                                        mgr26__std__lane24_strm0_data_valid  ;

  input                                         std__mgr26__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane24_strm1_data        ;
  output                                        mgr26__std__lane24_strm1_data_valid  ;

  input                                         std__mgr26__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane25_strm0_data        ;
  output                                        mgr26__std__lane25_strm0_data_valid  ;

  input                                         std__mgr26__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane25_strm1_data        ;
  output                                        mgr26__std__lane25_strm1_data_valid  ;

  input                                         std__mgr26__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane26_strm0_data        ;
  output                                        mgr26__std__lane26_strm0_data_valid  ;

  input                                         std__mgr26__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane26_strm1_data        ;
  output                                        mgr26__std__lane26_strm1_data_valid  ;

  input                                         std__mgr26__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane27_strm0_data        ;
  output                                        mgr26__std__lane27_strm0_data_valid  ;

  input                                         std__mgr26__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane27_strm1_data        ;
  output                                        mgr26__std__lane27_strm1_data_valid  ;

  input                                         std__mgr26__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane28_strm0_data        ;
  output                                        mgr26__std__lane28_strm0_data_valid  ;

  input                                         std__mgr26__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane28_strm1_data        ;
  output                                        mgr26__std__lane28_strm1_data_valid  ;

  input                                         std__mgr26__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane29_strm0_data        ;
  output                                        mgr26__std__lane29_strm0_data_valid  ;

  input                                         std__mgr26__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane29_strm1_data        ;
  output                                        mgr26__std__lane29_strm1_data_valid  ;

  input                                         std__mgr26__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane30_strm0_data        ;
  output                                        mgr26__std__lane30_strm0_data_valid  ;

  input                                         std__mgr26__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane30_strm1_data        ;
  output                                        mgr26__std__lane30_strm1_data_valid  ;

  input                                         std__mgr26__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane31_strm0_data        ;
  output                                        mgr26__std__lane31_strm0_data_valid  ;

  input                                         std__mgr26__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane31_strm1_data        ;
  output                                        mgr26__std__lane31_strm1_data_valid  ;

  input                                         std__mgr27__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane0_strm0_data        ;
  output                                        mgr27__std__lane0_strm0_data_valid  ;

  input                                         std__mgr27__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane0_strm1_data        ;
  output                                        mgr27__std__lane0_strm1_data_valid  ;

  input                                         std__mgr27__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane1_strm0_data        ;
  output                                        mgr27__std__lane1_strm0_data_valid  ;

  input                                         std__mgr27__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane1_strm1_data        ;
  output                                        mgr27__std__lane1_strm1_data_valid  ;

  input                                         std__mgr27__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane2_strm0_data        ;
  output                                        mgr27__std__lane2_strm0_data_valid  ;

  input                                         std__mgr27__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane2_strm1_data        ;
  output                                        mgr27__std__lane2_strm1_data_valid  ;

  input                                         std__mgr27__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane3_strm0_data        ;
  output                                        mgr27__std__lane3_strm0_data_valid  ;

  input                                         std__mgr27__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane3_strm1_data        ;
  output                                        mgr27__std__lane3_strm1_data_valid  ;

  input                                         std__mgr27__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane4_strm0_data        ;
  output                                        mgr27__std__lane4_strm0_data_valid  ;

  input                                         std__mgr27__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane4_strm1_data        ;
  output                                        mgr27__std__lane4_strm1_data_valid  ;

  input                                         std__mgr27__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane5_strm0_data        ;
  output                                        mgr27__std__lane5_strm0_data_valid  ;

  input                                         std__mgr27__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane5_strm1_data        ;
  output                                        mgr27__std__lane5_strm1_data_valid  ;

  input                                         std__mgr27__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane6_strm0_data        ;
  output                                        mgr27__std__lane6_strm0_data_valid  ;

  input                                         std__mgr27__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane6_strm1_data        ;
  output                                        mgr27__std__lane6_strm1_data_valid  ;

  input                                         std__mgr27__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane7_strm0_data        ;
  output                                        mgr27__std__lane7_strm0_data_valid  ;

  input                                         std__mgr27__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane7_strm1_data        ;
  output                                        mgr27__std__lane7_strm1_data_valid  ;

  input                                         std__mgr27__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane8_strm0_data        ;
  output                                        mgr27__std__lane8_strm0_data_valid  ;

  input                                         std__mgr27__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane8_strm1_data        ;
  output                                        mgr27__std__lane8_strm1_data_valid  ;

  input                                         std__mgr27__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane9_strm0_data        ;
  output                                        mgr27__std__lane9_strm0_data_valid  ;

  input                                         std__mgr27__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane9_strm1_data        ;
  output                                        mgr27__std__lane9_strm1_data_valid  ;

  input                                         std__mgr27__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane10_strm0_data        ;
  output                                        mgr27__std__lane10_strm0_data_valid  ;

  input                                         std__mgr27__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane10_strm1_data        ;
  output                                        mgr27__std__lane10_strm1_data_valid  ;

  input                                         std__mgr27__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane11_strm0_data        ;
  output                                        mgr27__std__lane11_strm0_data_valid  ;

  input                                         std__mgr27__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane11_strm1_data        ;
  output                                        mgr27__std__lane11_strm1_data_valid  ;

  input                                         std__mgr27__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane12_strm0_data        ;
  output                                        mgr27__std__lane12_strm0_data_valid  ;

  input                                         std__mgr27__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane12_strm1_data        ;
  output                                        mgr27__std__lane12_strm1_data_valid  ;

  input                                         std__mgr27__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane13_strm0_data        ;
  output                                        mgr27__std__lane13_strm0_data_valid  ;

  input                                         std__mgr27__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane13_strm1_data        ;
  output                                        mgr27__std__lane13_strm1_data_valid  ;

  input                                         std__mgr27__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane14_strm0_data        ;
  output                                        mgr27__std__lane14_strm0_data_valid  ;

  input                                         std__mgr27__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane14_strm1_data        ;
  output                                        mgr27__std__lane14_strm1_data_valid  ;

  input                                         std__mgr27__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane15_strm0_data        ;
  output                                        mgr27__std__lane15_strm0_data_valid  ;

  input                                         std__mgr27__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane15_strm1_data        ;
  output                                        mgr27__std__lane15_strm1_data_valid  ;

  input                                         std__mgr27__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane16_strm0_data        ;
  output                                        mgr27__std__lane16_strm0_data_valid  ;

  input                                         std__mgr27__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane16_strm1_data        ;
  output                                        mgr27__std__lane16_strm1_data_valid  ;

  input                                         std__mgr27__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane17_strm0_data        ;
  output                                        mgr27__std__lane17_strm0_data_valid  ;

  input                                         std__mgr27__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane17_strm1_data        ;
  output                                        mgr27__std__lane17_strm1_data_valid  ;

  input                                         std__mgr27__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane18_strm0_data        ;
  output                                        mgr27__std__lane18_strm0_data_valid  ;

  input                                         std__mgr27__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane18_strm1_data        ;
  output                                        mgr27__std__lane18_strm1_data_valid  ;

  input                                         std__mgr27__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane19_strm0_data        ;
  output                                        mgr27__std__lane19_strm0_data_valid  ;

  input                                         std__mgr27__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane19_strm1_data        ;
  output                                        mgr27__std__lane19_strm1_data_valid  ;

  input                                         std__mgr27__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane20_strm0_data        ;
  output                                        mgr27__std__lane20_strm0_data_valid  ;

  input                                         std__mgr27__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane20_strm1_data        ;
  output                                        mgr27__std__lane20_strm1_data_valid  ;

  input                                         std__mgr27__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane21_strm0_data        ;
  output                                        mgr27__std__lane21_strm0_data_valid  ;

  input                                         std__mgr27__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane21_strm1_data        ;
  output                                        mgr27__std__lane21_strm1_data_valid  ;

  input                                         std__mgr27__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane22_strm0_data        ;
  output                                        mgr27__std__lane22_strm0_data_valid  ;

  input                                         std__mgr27__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane22_strm1_data        ;
  output                                        mgr27__std__lane22_strm1_data_valid  ;

  input                                         std__mgr27__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane23_strm0_data        ;
  output                                        mgr27__std__lane23_strm0_data_valid  ;

  input                                         std__mgr27__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane23_strm1_data        ;
  output                                        mgr27__std__lane23_strm1_data_valid  ;

  input                                         std__mgr27__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane24_strm0_data        ;
  output                                        mgr27__std__lane24_strm0_data_valid  ;

  input                                         std__mgr27__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane24_strm1_data        ;
  output                                        mgr27__std__lane24_strm1_data_valid  ;

  input                                         std__mgr27__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane25_strm0_data        ;
  output                                        mgr27__std__lane25_strm0_data_valid  ;

  input                                         std__mgr27__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane25_strm1_data        ;
  output                                        mgr27__std__lane25_strm1_data_valid  ;

  input                                         std__mgr27__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane26_strm0_data        ;
  output                                        mgr27__std__lane26_strm0_data_valid  ;

  input                                         std__mgr27__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane26_strm1_data        ;
  output                                        mgr27__std__lane26_strm1_data_valid  ;

  input                                         std__mgr27__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane27_strm0_data        ;
  output                                        mgr27__std__lane27_strm0_data_valid  ;

  input                                         std__mgr27__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane27_strm1_data        ;
  output                                        mgr27__std__lane27_strm1_data_valid  ;

  input                                         std__mgr27__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane28_strm0_data        ;
  output                                        mgr27__std__lane28_strm0_data_valid  ;

  input                                         std__mgr27__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane28_strm1_data        ;
  output                                        mgr27__std__lane28_strm1_data_valid  ;

  input                                         std__mgr27__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane29_strm0_data        ;
  output                                        mgr27__std__lane29_strm0_data_valid  ;

  input                                         std__mgr27__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane29_strm1_data        ;
  output                                        mgr27__std__lane29_strm1_data_valid  ;

  input                                         std__mgr27__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane30_strm0_data        ;
  output                                        mgr27__std__lane30_strm0_data_valid  ;

  input                                         std__mgr27__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane30_strm1_data        ;
  output                                        mgr27__std__lane30_strm1_data_valid  ;

  input                                         std__mgr27__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane31_strm0_data        ;
  output                                        mgr27__std__lane31_strm0_data_valid  ;

  input                                         std__mgr27__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane31_strm1_data        ;
  output                                        mgr27__std__lane31_strm1_data_valid  ;

  input                                         std__mgr28__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane0_strm0_data        ;
  output                                        mgr28__std__lane0_strm0_data_valid  ;

  input                                         std__mgr28__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane0_strm1_data        ;
  output                                        mgr28__std__lane0_strm1_data_valid  ;

  input                                         std__mgr28__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane1_strm0_data        ;
  output                                        mgr28__std__lane1_strm0_data_valid  ;

  input                                         std__mgr28__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane1_strm1_data        ;
  output                                        mgr28__std__lane1_strm1_data_valid  ;

  input                                         std__mgr28__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane2_strm0_data        ;
  output                                        mgr28__std__lane2_strm0_data_valid  ;

  input                                         std__mgr28__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane2_strm1_data        ;
  output                                        mgr28__std__lane2_strm1_data_valid  ;

  input                                         std__mgr28__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane3_strm0_data        ;
  output                                        mgr28__std__lane3_strm0_data_valid  ;

  input                                         std__mgr28__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane3_strm1_data        ;
  output                                        mgr28__std__lane3_strm1_data_valid  ;

  input                                         std__mgr28__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane4_strm0_data        ;
  output                                        mgr28__std__lane4_strm0_data_valid  ;

  input                                         std__mgr28__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane4_strm1_data        ;
  output                                        mgr28__std__lane4_strm1_data_valid  ;

  input                                         std__mgr28__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane5_strm0_data        ;
  output                                        mgr28__std__lane5_strm0_data_valid  ;

  input                                         std__mgr28__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane5_strm1_data        ;
  output                                        mgr28__std__lane5_strm1_data_valid  ;

  input                                         std__mgr28__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane6_strm0_data        ;
  output                                        mgr28__std__lane6_strm0_data_valid  ;

  input                                         std__mgr28__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane6_strm1_data        ;
  output                                        mgr28__std__lane6_strm1_data_valid  ;

  input                                         std__mgr28__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane7_strm0_data        ;
  output                                        mgr28__std__lane7_strm0_data_valid  ;

  input                                         std__mgr28__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane7_strm1_data        ;
  output                                        mgr28__std__lane7_strm1_data_valid  ;

  input                                         std__mgr28__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane8_strm0_data        ;
  output                                        mgr28__std__lane8_strm0_data_valid  ;

  input                                         std__mgr28__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane8_strm1_data        ;
  output                                        mgr28__std__lane8_strm1_data_valid  ;

  input                                         std__mgr28__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane9_strm0_data        ;
  output                                        mgr28__std__lane9_strm0_data_valid  ;

  input                                         std__mgr28__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane9_strm1_data        ;
  output                                        mgr28__std__lane9_strm1_data_valid  ;

  input                                         std__mgr28__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane10_strm0_data        ;
  output                                        mgr28__std__lane10_strm0_data_valid  ;

  input                                         std__mgr28__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane10_strm1_data        ;
  output                                        mgr28__std__lane10_strm1_data_valid  ;

  input                                         std__mgr28__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane11_strm0_data        ;
  output                                        mgr28__std__lane11_strm0_data_valid  ;

  input                                         std__mgr28__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane11_strm1_data        ;
  output                                        mgr28__std__lane11_strm1_data_valid  ;

  input                                         std__mgr28__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane12_strm0_data        ;
  output                                        mgr28__std__lane12_strm0_data_valid  ;

  input                                         std__mgr28__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane12_strm1_data        ;
  output                                        mgr28__std__lane12_strm1_data_valid  ;

  input                                         std__mgr28__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane13_strm0_data        ;
  output                                        mgr28__std__lane13_strm0_data_valid  ;

  input                                         std__mgr28__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane13_strm1_data        ;
  output                                        mgr28__std__lane13_strm1_data_valid  ;

  input                                         std__mgr28__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane14_strm0_data        ;
  output                                        mgr28__std__lane14_strm0_data_valid  ;

  input                                         std__mgr28__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane14_strm1_data        ;
  output                                        mgr28__std__lane14_strm1_data_valid  ;

  input                                         std__mgr28__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane15_strm0_data        ;
  output                                        mgr28__std__lane15_strm0_data_valid  ;

  input                                         std__mgr28__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane15_strm1_data        ;
  output                                        mgr28__std__lane15_strm1_data_valid  ;

  input                                         std__mgr28__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane16_strm0_data        ;
  output                                        mgr28__std__lane16_strm0_data_valid  ;

  input                                         std__mgr28__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane16_strm1_data        ;
  output                                        mgr28__std__lane16_strm1_data_valid  ;

  input                                         std__mgr28__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane17_strm0_data        ;
  output                                        mgr28__std__lane17_strm0_data_valid  ;

  input                                         std__mgr28__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane17_strm1_data        ;
  output                                        mgr28__std__lane17_strm1_data_valid  ;

  input                                         std__mgr28__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane18_strm0_data        ;
  output                                        mgr28__std__lane18_strm0_data_valid  ;

  input                                         std__mgr28__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane18_strm1_data        ;
  output                                        mgr28__std__lane18_strm1_data_valid  ;

  input                                         std__mgr28__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane19_strm0_data        ;
  output                                        mgr28__std__lane19_strm0_data_valid  ;

  input                                         std__mgr28__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane19_strm1_data        ;
  output                                        mgr28__std__lane19_strm1_data_valid  ;

  input                                         std__mgr28__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane20_strm0_data        ;
  output                                        mgr28__std__lane20_strm0_data_valid  ;

  input                                         std__mgr28__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane20_strm1_data        ;
  output                                        mgr28__std__lane20_strm1_data_valid  ;

  input                                         std__mgr28__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane21_strm0_data        ;
  output                                        mgr28__std__lane21_strm0_data_valid  ;

  input                                         std__mgr28__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane21_strm1_data        ;
  output                                        mgr28__std__lane21_strm1_data_valid  ;

  input                                         std__mgr28__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane22_strm0_data        ;
  output                                        mgr28__std__lane22_strm0_data_valid  ;

  input                                         std__mgr28__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane22_strm1_data        ;
  output                                        mgr28__std__lane22_strm1_data_valid  ;

  input                                         std__mgr28__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane23_strm0_data        ;
  output                                        mgr28__std__lane23_strm0_data_valid  ;

  input                                         std__mgr28__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane23_strm1_data        ;
  output                                        mgr28__std__lane23_strm1_data_valid  ;

  input                                         std__mgr28__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane24_strm0_data        ;
  output                                        mgr28__std__lane24_strm0_data_valid  ;

  input                                         std__mgr28__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane24_strm1_data        ;
  output                                        mgr28__std__lane24_strm1_data_valid  ;

  input                                         std__mgr28__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane25_strm0_data        ;
  output                                        mgr28__std__lane25_strm0_data_valid  ;

  input                                         std__mgr28__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane25_strm1_data        ;
  output                                        mgr28__std__lane25_strm1_data_valid  ;

  input                                         std__mgr28__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane26_strm0_data        ;
  output                                        mgr28__std__lane26_strm0_data_valid  ;

  input                                         std__mgr28__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane26_strm1_data        ;
  output                                        mgr28__std__lane26_strm1_data_valid  ;

  input                                         std__mgr28__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane27_strm0_data        ;
  output                                        mgr28__std__lane27_strm0_data_valid  ;

  input                                         std__mgr28__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane27_strm1_data        ;
  output                                        mgr28__std__lane27_strm1_data_valid  ;

  input                                         std__mgr28__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane28_strm0_data        ;
  output                                        mgr28__std__lane28_strm0_data_valid  ;

  input                                         std__mgr28__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane28_strm1_data        ;
  output                                        mgr28__std__lane28_strm1_data_valid  ;

  input                                         std__mgr28__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane29_strm0_data        ;
  output                                        mgr28__std__lane29_strm0_data_valid  ;

  input                                         std__mgr28__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane29_strm1_data        ;
  output                                        mgr28__std__lane29_strm1_data_valid  ;

  input                                         std__mgr28__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane30_strm0_data        ;
  output                                        mgr28__std__lane30_strm0_data_valid  ;

  input                                         std__mgr28__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane30_strm1_data        ;
  output                                        mgr28__std__lane30_strm1_data_valid  ;

  input                                         std__mgr28__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane31_strm0_data        ;
  output                                        mgr28__std__lane31_strm0_data_valid  ;

  input                                         std__mgr28__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane31_strm1_data        ;
  output                                        mgr28__std__lane31_strm1_data_valid  ;

  input                                         std__mgr29__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane0_strm0_data        ;
  output                                        mgr29__std__lane0_strm0_data_valid  ;

  input                                         std__mgr29__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane0_strm1_data        ;
  output                                        mgr29__std__lane0_strm1_data_valid  ;

  input                                         std__mgr29__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane1_strm0_data        ;
  output                                        mgr29__std__lane1_strm0_data_valid  ;

  input                                         std__mgr29__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane1_strm1_data        ;
  output                                        mgr29__std__lane1_strm1_data_valid  ;

  input                                         std__mgr29__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane2_strm0_data        ;
  output                                        mgr29__std__lane2_strm0_data_valid  ;

  input                                         std__mgr29__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane2_strm1_data        ;
  output                                        mgr29__std__lane2_strm1_data_valid  ;

  input                                         std__mgr29__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane3_strm0_data        ;
  output                                        mgr29__std__lane3_strm0_data_valid  ;

  input                                         std__mgr29__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane3_strm1_data        ;
  output                                        mgr29__std__lane3_strm1_data_valid  ;

  input                                         std__mgr29__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane4_strm0_data        ;
  output                                        mgr29__std__lane4_strm0_data_valid  ;

  input                                         std__mgr29__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane4_strm1_data        ;
  output                                        mgr29__std__lane4_strm1_data_valid  ;

  input                                         std__mgr29__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane5_strm0_data        ;
  output                                        mgr29__std__lane5_strm0_data_valid  ;

  input                                         std__mgr29__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane5_strm1_data        ;
  output                                        mgr29__std__lane5_strm1_data_valid  ;

  input                                         std__mgr29__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane6_strm0_data        ;
  output                                        mgr29__std__lane6_strm0_data_valid  ;

  input                                         std__mgr29__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane6_strm1_data        ;
  output                                        mgr29__std__lane6_strm1_data_valid  ;

  input                                         std__mgr29__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane7_strm0_data        ;
  output                                        mgr29__std__lane7_strm0_data_valid  ;

  input                                         std__mgr29__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane7_strm1_data        ;
  output                                        mgr29__std__lane7_strm1_data_valid  ;

  input                                         std__mgr29__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane8_strm0_data        ;
  output                                        mgr29__std__lane8_strm0_data_valid  ;

  input                                         std__mgr29__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane8_strm1_data        ;
  output                                        mgr29__std__lane8_strm1_data_valid  ;

  input                                         std__mgr29__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane9_strm0_data        ;
  output                                        mgr29__std__lane9_strm0_data_valid  ;

  input                                         std__mgr29__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane9_strm1_data        ;
  output                                        mgr29__std__lane9_strm1_data_valid  ;

  input                                         std__mgr29__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane10_strm0_data        ;
  output                                        mgr29__std__lane10_strm0_data_valid  ;

  input                                         std__mgr29__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane10_strm1_data        ;
  output                                        mgr29__std__lane10_strm1_data_valid  ;

  input                                         std__mgr29__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane11_strm0_data        ;
  output                                        mgr29__std__lane11_strm0_data_valid  ;

  input                                         std__mgr29__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane11_strm1_data        ;
  output                                        mgr29__std__lane11_strm1_data_valid  ;

  input                                         std__mgr29__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane12_strm0_data        ;
  output                                        mgr29__std__lane12_strm0_data_valid  ;

  input                                         std__mgr29__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane12_strm1_data        ;
  output                                        mgr29__std__lane12_strm1_data_valid  ;

  input                                         std__mgr29__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane13_strm0_data        ;
  output                                        mgr29__std__lane13_strm0_data_valid  ;

  input                                         std__mgr29__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane13_strm1_data        ;
  output                                        mgr29__std__lane13_strm1_data_valid  ;

  input                                         std__mgr29__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane14_strm0_data        ;
  output                                        mgr29__std__lane14_strm0_data_valid  ;

  input                                         std__mgr29__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane14_strm1_data        ;
  output                                        mgr29__std__lane14_strm1_data_valid  ;

  input                                         std__mgr29__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane15_strm0_data        ;
  output                                        mgr29__std__lane15_strm0_data_valid  ;

  input                                         std__mgr29__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane15_strm1_data        ;
  output                                        mgr29__std__lane15_strm1_data_valid  ;

  input                                         std__mgr29__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane16_strm0_data        ;
  output                                        mgr29__std__lane16_strm0_data_valid  ;

  input                                         std__mgr29__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane16_strm1_data        ;
  output                                        mgr29__std__lane16_strm1_data_valid  ;

  input                                         std__mgr29__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane17_strm0_data        ;
  output                                        mgr29__std__lane17_strm0_data_valid  ;

  input                                         std__mgr29__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane17_strm1_data        ;
  output                                        mgr29__std__lane17_strm1_data_valid  ;

  input                                         std__mgr29__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane18_strm0_data        ;
  output                                        mgr29__std__lane18_strm0_data_valid  ;

  input                                         std__mgr29__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane18_strm1_data        ;
  output                                        mgr29__std__lane18_strm1_data_valid  ;

  input                                         std__mgr29__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane19_strm0_data        ;
  output                                        mgr29__std__lane19_strm0_data_valid  ;

  input                                         std__mgr29__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane19_strm1_data        ;
  output                                        mgr29__std__lane19_strm1_data_valid  ;

  input                                         std__mgr29__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane20_strm0_data        ;
  output                                        mgr29__std__lane20_strm0_data_valid  ;

  input                                         std__mgr29__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane20_strm1_data        ;
  output                                        mgr29__std__lane20_strm1_data_valid  ;

  input                                         std__mgr29__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane21_strm0_data        ;
  output                                        mgr29__std__lane21_strm0_data_valid  ;

  input                                         std__mgr29__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane21_strm1_data        ;
  output                                        mgr29__std__lane21_strm1_data_valid  ;

  input                                         std__mgr29__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane22_strm0_data        ;
  output                                        mgr29__std__lane22_strm0_data_valid  ;

  input                                         std__mgr29__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane22_strm1_data        ;
  output                                        mgr29__std__lane22_strm1_data_valid  ;

  input                                         std__mgr29__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane23_strm0_data        ;
  output                                        mgr29__std__lane23_strm0_data_valid  ;

  input                                         std__mgr29__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane23_strm1_data        ;
  output                                        mgr29__std__lane23_strm1_data_valid  ;

  input                                         std__mgr29__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane24_strm0_data        ;
  output                                        mgr29__std__lane24_strm0_data_valid  ;

  input                                         std__mgr29__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane24_strm1_data        ;
  output                                        mgr29__std__lane24_strm1_data_valid  ;

  input                                         std__mgr29__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane25_strm0_data        ;
  output                                        mgr29__std__lane25_strm0_data_valid  ;

  input                                         std__mgr29__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane25_strm1_data        ;
  output                                        mgr29__std__lane25_strm1_data_valid  ;

  input                                         std__mgr29__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane26_strm0_data        ;
  output                                        mgr29__std__lane26_strm0_data_valid  ;

  input                                         std__mgr29__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane26_strm1_data        ;
  output                                        mgr29__std__lane26_strm1_data_valid  ;

  input                                         std__mgr29__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane27_strm0_data        ;
  output                                        mgr29__std__lane27_strm0_data_valid  ;

  input                                         std__mgr29__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane27_strm1_data        ;
  output                                        mgr29__std__lane27_strm1_data_valid  ;

  input                                         std__mgr29__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane28_strm0_data        ;
  output                                        mgr29__std__lane28_strm0_data_valid  ;

  input                                         std__mgr29__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane28_strm1_data        ;
  output                                        mgr29__std__lane28_strm1_data_valid  ;

  input                                         std__mgr29__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane29_strm0_data        ;
  output                                        mgr29__std__lane29_strm0_data_valid  ;

  input                                         std__mgr29__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane29_strm1_data        ;
  output                                        mgr29__std__lane29_strm1_data_valid  ;

  input                                         std__mgr29__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane30_strm0_data        ;
  output                                        mgr29__std__lane30_strm0_data_valid  ;

  input                                         std__mgr29__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane30_strm1_data        ;
  output                                        mgr29__std__lane30_strm1_data_valid  ;

  input                                         std__mgr29__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane31_strm0_data        ;
  output                                        mgr29__std__lane31_strm0_data_valid  ;

  input                                         std__mgr29__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane31_strm1_data        ;
  output                                        mgr29__std__lane31_strm1_data_valid  ;

  input                                         std__mgr30__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane0_strm0_data        ;
  output                                        mgr30__std__lane0_strm0_data_valid  ;

  input                                         std__mgr30__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane0_strm1_data        ;
  output                                        mgr30__std__lane0_strm1_data_valid  ;

  input                                         std__mgr30__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane1_strm0_data        ;
  output                                        mgr30__std__lane1_strm0_data_valid  ;

  input                                         std__mgr30__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane1_strm1_data        ;
  output                                        mgr30__std__lane1_strm1_data_valid  ;

  input                                         std__mgr30__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane2_strm0_data        ;
  output                                        mgr30__std__lane2_strm0_data_valid  ;

  input                                         std__mgr30__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane2_strm1_data        ;
  output                                        mgr30__std__lane2_strm1_data_valid  ;

  input                                         std__mgr30__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane3_strm0_data        ;
  output                                        mgr30__std__lane3_strm0_data_valid  ;

  input                                         std__mgr30__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane3_strm1_data        ;
  output                                        mgr30__std__lane3_strm1_data_valid  ;

  input                                         std__mgr30__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane4_strm0_data        ;
  output                                        mgr30__std__lane4_strm0_data_valid  ;

  input                                         std__mgr30__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane4_strm1_data        ;
  output                                        mgr30__std__lane4_strm1_data_valid  ;

  input                                         std__mgr30__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane5_strm0_data        ;
  output                                        mgr30__std__lane5_strm0_data_valid  ;

  input                                         std__mgr30__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane5_strm1_data        ;
  output                                        mgr30__std__lane5_strm1_data_valid  ;

  input                                         std__mgr30__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane6_strm0_data        ;
  output                                        mgr30__std__lane6_strm0_data_valid  ;

  input                                         std__mgr30__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane6_strm1_data        ;
  output                                        mgr30__std__lane6_strm1_data_valid  ;

  input                                         std__mgr30__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane7_strm0_data        ;
  output                                        mgr30__std__lane7_strm0_data_valid  ;

  input                                         std__mgr30__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane7_strm1_data        ;
  output                                        mgr30__std__lane7_strm1_data_valid  ;

  input                                         std__mgr30__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane8_strm0_data        ;
  output                                        mgr30__std__lane8_strm0_data_valid  ;

  input                                         std__mgr30__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane8_strm1_data        ;
  output                                        mgr30__std__lane8_strm1_data_valid  ;

  input                                         std__mgr30__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane9_strm0_data        ;
  output                                        mgr30__std__lane9_strm0_data_valid  ;

  input                                         std__mgr30__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane9_strm1_data        ;
  output                                        mgr30__std__lane9_strm1_data_valid  ;

  input                                         std__mgr30__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane10_strm0_data        ;
  output                                        mgr30__std__lane10_strm0_data_valid  ;

  input                                         std__mgr30__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane10_strm1_data        ;
  output                                        mgr30__std__lane10_strm1_data_valid  ;

  input                                         std__mgr30__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane11_strm0_data        ;
  output                                        mgr30__std__lane11_strm0_data_valid  ;

  input                                         std__mgr30__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane11_strm1_data        ;
  output                                        mgr30__std__lane11_strm1_data_valid  ;

  input                                         std__mgr30__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane12_strm0_data        ;
  output                                        mgr30__std__lane12_strm0_data_valid  ;

  input                                         std__mgr30__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane12_strm1_data        ;
  output                                        mgr30__std__lane12_strm1_data_valid  ;

  input                                         std__mgr30__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane13_strm0_data        ;
  output                                        mgr30__std__lane13_strm0_data_valid  ;

  input                                         std__mgr30__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane13_strm1_data        ;
  output                                        mgr30__std__lane13_strm1_data_valid  ;

  input                                         std__mgr30__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane14_strm0_data        ;
  output                                        mgr30__std__lane14_strm0_data_valid  ;

  input                                         std__mgr30__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane14_strm1_data        ;
  output                                        mgr30__std__lane14_strm1_data_valid  ;

  input                                         std__mgr30__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane15_strm0_data        ;
  output                                        mgr30__std__lane15_strm0_data_valid  ;

  input                                         std__mgr30__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane15_strm1_data        ;
  output                                        mgr30__std__lane15_strm1_data_valid  ;

  input                                         std__mgr30__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane16_strm0_data        ;
  output                                        mgr30__std__lane16_strm0_data_valid  ;

  input                                         std__mgr30__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane16_strm1_data        ;
  output                                        mgr30__std__lane16_strm1_data_valid  ;

  input                                         std__mgr30__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane17_strm0_data        ;
  output                                        mgr30__std__lane17_strm0_data_valid  ;

  input                                         std__mgr30__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane17_strm1_data        ;
  output                                        mgr30__std__lane17_strm1_data_valid  ;

  input                                         std__mgr30__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane18_strm0_data        ;
  output                                        mgr30__std__lane18_strm0_data_valid  ;

  input                                         std__mgr30__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane18_strm1_data        ;
  output                                        mgr30__std__lane18_strm1_data_valid  ;

  input                                         std__mgr30__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane19_strm0_data        ;
  output                                        mgr30__std__lane19_strm0_data_valid  ;

  input                                         std__mgr30__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane19_strm1_data        ;
  output                                        mgr30__std__lane19_strm1_data_valid  ;

  input                                         std__mgr30__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane20_strm0_data        ;
  output                                        mgr30__std__lane20_strm0_data_valid  ;

  input                                         std__mgr30__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane20_strm1_data        ;
  output                                        mgr30__std__lane20_strm1_data_valid  ;

  input                                         std__mgr30__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane21_strm0_data        ;
  output                                        mgr30__std__lane21_strm0_data_valid  ;

  input                                         std__mgr30__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane21_strm1_data        ;
  output                                        mgr30__std__lane21_strm1_data_valid  ;

  input                                         std__mgr30__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane22_strm0_data        ;
  output                                        mgr30__std__lane22_strm0_data_valid  ;

  input                                         std__mgr30__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane22_strm1_data        ;
  output                                        mgr30__std__lane22_strm1_data_valid  ;

  input                                         std__mgr30__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane23_strm0_data        ;
  output                                        mgr30__std__lane23_strm0_data_valid  ;

  input                                         std__mgr30__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane23_strm1_data        ;
  output                                        mgr30__std__lane23_strm1_data_valid  ;

  input                                         std__mgr30__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane24_strm0_data        ;
  output                                        mgr30__std__lane24_strm0_data_valid  ;

  input                                         std__mgr30__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane24_strm1_data        ;
  output                                        mgr30__std__lane24_strm1_data_valid  ;

  input                                         std__mgr30__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane25_strm0_data        ;
  output                                        mgr30__std__lane25_strm0_data_valid  ;

  input                                         std__mgr30__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane25_strm1_data        ;
  output                                        mgr30__std__lane25_strm1_data_valid  ;

  input                                         std__mgr30__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane26_strm0_data        ;
  output                                        mgr30__std__lane26_strm0_data_valid  ;

  input                                         std__mgr30__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane26_strm1_data        ;
  output                                        mgr30__std__lane26_strm1_data_valid  ;

  input                                         std__mgr30__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane27_strm0_data        ;
  output                                        mgr30__std__lane27_strm0_data_valid  ;

  input                                         std__mgr30__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane27_strm1_data        ;
  output                                        mgr30__std__lane27_strm1_data_valid  ;

  input                                         std__mgr30__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane28_strm0_data        ;
  output                                        mgr30__std__lane28_strm0_data_valid  ;

  input                                         std__mgr30__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane28_strm1_data        ;
  output                                        mgr30__std__lane28_strm1_data_valid  ;

  input                                         std__mgr30__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane29_strm0_data        ;
  output                                        mgr30__std__lane29_strm0_data_valid  ;

  input                                         std__mgr30__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane29_strm1_data        ;
  output                                        mgr30__std__lane29_strm1_data_valid  ;

  input                                         std__mgr30__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane30_strm0_data        ;
  output                                        mgr30__std__lane30_strm0_data_valid  ;

  input                                         std__mgr30__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane30_strm1_data        ;
  output                                        mgr30__std__lane30_strm1_data_valid  ;

  input                                         std__mgr30__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane31_strm0_data        ;
  output                                        mgr30__std__lane31_strm0_data_valid  ;

  input                                         std__mgr30__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane31_strm1_data        ;
  output                                        mgr30__std__lane31_strm1_data_valid  ;

  input                                         std__mgr31__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane0_strm0_data        ;
  output                                        mgr31__std__lane0_strm0_data_valid  ;

  input                                         std__mgr31__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane0_strm1_data        ;
  output                                        mgr31__std__lane0_strm1_data_valid  ;

  input                                         std__mgr31__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane1_strm0_data        ;
  output                                        mgr31__std__lane1_strm0_data_valid  ;

  input                                         std__mgr31__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane1_strm1_data        ;
  output                                        mgr31__std__lane1_strm1_data_valid  ;

  input                                         std__mgr31__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane2_strm0_data        ;
  output                                        mgr31__std__lane2_strm0_data_valid  ;

  input                                         std__mgr31__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane2_strm1_data        ;
  output                                        mgr31__std__lane2_strm1_data_valid  ;

  input                                         std__mgr31__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane3_strm0_data        ;
  output                                        mgr31__std__lane3_strm0_data_valid  ;

  input                                         std__mgr31__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane3_strm1_data        ;
  output                                        mgr31__std__lane3_strm1_data_valid  ;

  input                                         std__mgr31__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane4_strm0_data        ;
  output                                        mgr31__std__lane4_strm0_data_valid  ;

  input                                         std__mgr31__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane4_strm1_data        ;
  output                                        mgr31__std__lane4_strm1_data_valid  ;

  input                                         std__mgr31__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane5_strm0_data        ;
  output                                        mgr31__std__lane5_strm0_data_valid  ;

  input                                         std__mgr31__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane5_strm1_data        ;
  output                                        mgr31__std__lane5_strm1_data_valid  ;

  input                                         std__mgr31__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane6_strm0_data        ;
  output                                        mgr31__std__lane6_strm0_data_valid  ;

  input                                         std__mgr31__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane6_strm1_data        ;
  output                                        mgr31__std__lane6_strm1_data_valid  ;

  input                                         std__mgr31__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane7_strm0_data        ;
  output                                        mgr31__std__lane7_strm0_data_valid  ;

  input                                         std__mgr31__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane7_strm1_data        ;
  output                                        mgr31__std__lane7_strm1_data_valid  ;

  input                                         std__mgr31__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane8_strm0_data        ;
  output                                        mgr31__std__lane8_strm0_data_valid  ;

  input                                         std__mgr31__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane8_strm1_data        ;
  output                                        mgr31__std__lane8_strm1_data_valid  ;

  input                                         std__mgr31__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane9_strm0_data        ;
  output                                        mgr31__std__lane9_strm0_data_valid  ;

  input                                         std__mgr31__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane9_strm1_data        ;
  output                                        mgr31__std__lane9_strm1_data_valid  ;

  input                                         std__mgr31__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane10_strm0_data        ;
  output                                        mgr31__std__lane10_strm0_data_valid  ;

  input                                         std__mgr31__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane10_strm1_data        ;
  output                                        mgr31__std__lane10_strm1_data_valid  ;

  input                                         std__mgr31__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane11_strm0_data        ;
  output                                        mgr31__std__lane11_strm0_data_valid  ;

  input                                         std__mgr31__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane11_strm1_data        ;
  output                                        mgr31__std__lane11_strm1_data_valid  ;

  input                                         std__mgr31__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane12_strm0_data        ;
  output                                        mgr31__std__lane12_strm0_data_valid  ;

  input                                         std__mgr31__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane12_strm1_data        ;
  output                                        mgr31__std__lane12_strm1_data_valid  ;

  input                                         std__mgr31__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane13_strm0_data        ;
  output                                        mgr31__std__lane13_strm0_data_valid  ;

  input                                         std__mgr31__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane13_strm1_data        ;
  output                                        mgr31__std__lane13_strm1_data_valid  ;

  input                                         std__mgr31__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane14_strm0_data        ;
  output                                        mgr31__std__lane14_strm0_data_valid  ;

  input                                         std__mgr31__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane14_strm1_data        ;
  output                                        mgr31__std__lane14_strm1_data_valid  ;

  input                                         std__mgr31__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane15_strm0_data        ;
  output                                        mgr31__std__lane15_strm0_data_valid  ;

  input                                         std__mgr31__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane15_strm1_data        ;
  output                                        mgr31__std__lane15_strm1_data_valid  ;

  input                                         std__mgr31__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane16_strm0_data        ;
  output                                        mgr31__std__lane16_strm0_data_valid  ;

  input                                         std__mgr31__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane16_strm1_data        ;
  output                                        mgr31__std__lane16_strm1_data_valid  ;

  input                                         std__mgr31__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane17_strm0_data        ;
  output                                        mgr31__std__lane17_strm0_data_valid  ;

  input                                         std__mgr31__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane17_strm1_data        ;
  output                                        mgr31__std__lane17_strm1_data_valid  ;

  input                                         std__mgr31__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane18_strm0_data        ;
  output                                        mgr31__std__lane18_strm0_data_valid  ;

  input                                         std__mgr31__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane18_strm1_data        ;
  output                                        mgr31__std__lane18_strm1_data_valid  ;

  input                                         std__mgr31__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane19_strm0_data        ;
  output                                        mgr31__std__lane19_strm0_data_valid  ;

  input                                         std__mgr31__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane19_strm1_data        ;
  output                                        mgr31__std__lane19_strm1_data_valid  ;

  input                                         std__mgr31__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane20_strm0_data        ;
  output                                        mgr31__std__lane20_strm0_data_valid  ;

  input                                         std__mgr31__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane20_strm1_data        ;
  output                                        mgr31__std__lane20_strm1_data_valid  ;

  input                                         std__mgr31__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane21_strm0_data        ;
  output                                        mgr31__std__lane21_strm0_data_valid  ;

  input                                         std__mgr31__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane21_strm1_data        ;
  output                                        mgr31__std__lane21_strm1_data_valid  ;

  input                                         std__mgr31__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane22_strm0_data        ;
  output                                        mgr31__std__lane22_strm0_data_valid  ;

  input                                         std__mgr31__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane22_strm1_data        ;
  output                                        mgr31__std__lane22_strm1_data_valid  ;

  input                                         std__mgr31__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane23_strm0_data        ;
  output                                        mgr31__std__lane23_strm0_data_valid  ;

  input                                         std__mgr31__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane23_strm1_data        ;
  output                                        mgr31__std__lane23_strm1_data_valid  ;

  input                                         std__mgr31__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane24_strm0_data        ;
  output                                        mgr31__std__lane24_strm0_data_valid  ;

  input                                         std__mgr31__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane24_strm1_data        ;
  output                                        mgr31__std__lane24_strm1_data_valid  ;

  input                                         std__mgr31__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane25_strm0_data        ;
  output                                        mgr31__std__lane25_strm0_data_valid  ;

  input                                         std__mgr31__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane25_strm1_data        ;
  output                                        mgr31__std__lane25_strm1_data_valid  ;

  input                                         std__mgr31__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane26_strm0_data        ;
  output                                        mgr31__std__lane26_strm0_data_valid  ;

  input                                         std__mgr31__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane26_strm1_data        ;
  output                                        mgr31__std__lane26_strm1_data_valid  ;

  input                                         std__mgr31__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane27_strm0_data        ;
  output                                        mgr31__std__lane27_strm0_data_valid  ;

  input                                         std__mgr31__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane27_strm1_data        ;
  output                                        mgr31__std__lane27_strm1_data_valid  ;

  input                                         std__mgr31__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane28_strm0_data        ;
  output                                        mgr31__std__lane28_strm0_data_valid  ;

  input                                         std__mgr31__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane28_strm1_data        ;
  output                                        mgr31__std__lane28_strm1_data_valid  ;

  input                                         std__mgr31__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane29_strm0_data        ;
  output                                        mgr31__std__lane29_strm0_data_valid  ;

  input                                         std__mgr31__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane29_strm1_data        ;
  output                                        mgr31__std__lane29_strm1_data_valid  ;

  input                                         std__mgr31__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane30_strm0_data        ;
  output                                        mgr31__std__lane30_strm0_data_valid  ;

  input                                         std__mgr31__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane30_strm1_data        ;
  output                                        mgr31__std__lane30_strm1_data_valid  ;

  input                                         std__mgr31__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane31_strm0_data        ;
  output                                        mgr31__std__lane31_strm0_data_valid  ;

  input                                         std__mgr31__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane31_strm1_data        ;
  output                                        mgr31__std__lane31_strm1_data_valid  ;

  input                                         std__mgr32__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane0_strm0_data        ;
  output                                        mgr32__std__lane0_strm0_data_valid  ;

  input                                         std__mgr32__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane0_strm1_data        ;
  output                                        mgr32__std__lane0_strm1_data_valid  ;

  input                                         std__mgr32__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane1_strm0_data        ;
  output                                        mgr32__std__lane1_strm0_data_valid  ;

  input                                         std__mgr32__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane1_strm1_data        ;
  output                                        mgr32__std__lane1_strm1_data_valid  ;

  input                                         std__mgr32__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane2_strm0_data        ;
  output                                        mgr32__std__lane2_strm0_data_valid  ;

  input                                         std__mgr32__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane2_strm1_data        ;
  output                                        mgr32__std__lane2_strm1_data_valid  ;

  input                                         std__mgr32__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane3_strm0_data        ;
  output                                        mgr32__std__lane3_strm0_data_valid  ;

  input                                         std__mgr32__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane3_strm1_data        ;
  output                                        mgr32__std__lane3_strm1_data_valid  ;

  input                                         std__mgr32__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane4_strm0_data        ;
  output                                        mgr32__std__lane4_strm0_data_valid  ;

  input                                         std__mgr32__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane4_strm1_data        ;
  output                                        mgr32__std__lane4_strm1_data_valid  ;

  input                                         std__mgr32__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane5_strm0_data        ;
  output                                        mgr32__std__lane5_strm0_data_valid  ;

  input                                         std__mgr32__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane5_strm1_data        ;
  output                                        mgr32__std__lane5_strm1_data_valid  ;

  input                                         std__mgr32__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane6_strm0_data        ;
  output                                        mgr32__std__lane6_strm0_data_valid  ;

  input                                         std__mgr32__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane6_strm1_data        ;
  output                                        mgr32__std__lane6_strm1_data_valid  ;

  input                                         std__mgr32__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane7_strm0_data        ;
  output                                        mgr32__std__lane7_strm0_data_valid  ;

  input                                         std__mgr32__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane7_strm1_data        ;
  output                                        mgr32__std__lane7_strm1_data_valid  ;

  input                                         std__mgr32__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane8_strm0_data        ;
  output                                        mgr32__std__lane8_strm0_data_valid  ;

  input                                         std__mgr32__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane8_strm1_data        ;
  output                                        mgr32__std__lane8_strm1_data_valid  ;

  input                                         std__mgr32__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane9_strm0_data        ;
  output                                        mgr32__std__lane9_strm0_data_valid  ;

  input                                         std__mgr32__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane9_strm1_data        ;
  output                                        mgr32__std__lane9_strm1_data_valid  ;

  input                                         std__mgr32__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane10_strm0_data        ;
  output                                        mgr32__std__lane10_strm0_data_valid  ;

  input                                         std__mgr32__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane10_strm1_data        ;
  output                                        mgr32__std__lane10_strm1_data_valid  ;

  input                                         std__mgr32__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane11_strm0_data        ;
  output                                        mgr32__std__lane11_strm0_data_valid  ;

  input                                         std__mgr32__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane11_strm1_data        ;
  output                                        mgr32__std__lane11_strm1_data_valid  ;

  input                                         std__mgr32__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane12_strm0_data        ;
  output                                        mgr32__std__lane12_strm0_data_valid  ;

  input                                         std__mgr32__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane12_strm1_data        ;
  output                                        mgr32__std__lane12_strm1_data_valid  ;

  input                                         std__mgr32__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane13_strm0_data        ;
  output                                        mgr32__std__lane13_strm0_data_valid  ;

  input                                         std__mgr32__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane13_strm1_data        ;
  output                                        mgr32__std__lane13_strm1_data_valid  ;

  input                                         std__mgr32__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane14_strm0_data        ;
  output                                        mgr32__std__lane14_strm0_data_valid  ;

  input                                         std__mgr32__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane14_strm1_data        ;
  output                                        mgr32__std__lane14_strm1_data_valid  ;

  input                                         std__mgr32__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane15_strm0_data        ;
  output                                        mgr32__std__lane15_strm0_data_valid  ;

  input                                         std__mgr32__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane15_strm1_data        ;
  output                                        mgr32__std__lane15_strm1_data_valid  ;

  input                                         std__mgr32__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane16_strm0_data        ;
  output                                        mgr32__std__lane16_strm0_data_valid  ;

  input                                         std__mgr32__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane16_strm1_data        ;
  output                                        mgr32__std__lane16_strm1_data_valid  ;

  input                                         std__mgr32__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane17_strm0_data        ;
  output                                        mgr32__std__lane17_strm0_data_valid  ;

  input                                         std__mgr32__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane17_strm1_data        ;
  output                                        mgr32__std__lane17_strm1_data_valid  ;

  input                                         std__mgr32__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane18_strm0_data        ;
  output                                        mgr32__std__lane18_strm0_data_valid  ;

  input                                         std__mgr32__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane18_strm1_data        ;
  output                                        mgr32__std__lane18_strm1_data_valid  ;

  input                                         std__mgr32__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane19_strm0_data        ;
  output                                        mgr32__std__lane19_strm0_data_valid  ;

  input                                         std__mgr32__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane19_strm1_data        ;
  output                                        mgr32__std__lane19_strm1_data_valid  ;

  input                                         std__mgr32__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane20_strm0_data        ;
  output                                        mgr32__std__lane20_strm0_data_valid  ;

  input                                         std__mgr32__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane20_strm1_data        ;
  output                                        mgr32__std__lane20_strm1_data_valid  ;

  input                                         std__mgr32__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane21_strm0_data        ;
  output                                        mgr32__std__lane21_strm0_data_valid  ;

  input                                         std__mgr32__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane21_strm1_data        ;
  output                                        mgr32__std__lane21_strm1_data_valid  ;

  input                                         std__mgr32__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane22_strm0_data        ;
  output                                        mgr32__std__lane22_strm0_data_valid  ;

  input                                         std__mgr32__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane22_strm1_data        ;
  output                                        mgr32__std__lane22_strm1_data_valid  ;

  input                                         std__mgr32__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane23_strm0_data        ;
  output                                        mgr32__std__lane23_strm0_data_valid  ;

  input                                         std__mgr32__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane23_strm1_data        ;
  output                                        mgr32__std__lane23_strm1_data_valid  ;

  input                                         std__mgr32__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane24_strm0_data        ;
  output                                        mgr32__std__lane24_strm0_data_valid  ;

  input                                         std__mgr32__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane24_strm1_data        ;
  output                                        mgr32__std__lane24_strm1_data_valid  ;

  input                                         std__mgr32__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane25_strm0_data        ;
  output                                        mgr32__std__lane25_strm0_data_valid  ;

  input                                         std__mgr32__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane25_strm1_data        ;
  output                                        mgr32__std__lane25_strm1_data_valid  ;

  input                                         std__mgr32__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane26_strm0_data        ;
  output                                        mgr32__std__lane26_strm0_data_valid  ;

  input                                         std__mgr32__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane26_strm1_data        ;
  output                                        mgr32__std__lane26_strm1_data_valid  ;

  input                                         std__mgr32__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane27_strm0_data        ;
  output                                        mgr32__std__lane27_strm0_data_valid  ;

  input                                         std__mgr32__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane27_strm1_data        ;
  output                                        mgr32__std__lane27_strm1_data_valid  ;

  input                                         std__mgr32__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane28_strm0_data        ;
  output                                        mgr32__std__lane28_strm0_data_valid  ;

  input                                         std__mgr32__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane28_strm1_data        ;
  output                                        mgr32__std__lane28_strm1_data_valid  ;

  input                                         std__mgr32__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane29_strm0_data        ;
  output                                        mgr32__std__lane29_strm0_data_valid  ;

  input                                         std__mgr32__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane29_strm1_data        ;
  output                                        mgr32__std__lane29_strm1_data_valid  ;

  input                                         std__mgr32__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane30_strm0_data        ;
  output                                        mgr32__std__lane30_strm0_data_valid  ;

  input                                         std__mgr32__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane30_strm1_data        ;
  output                                        mgr32__std__lane30_strm1_data_valid  ;

  input                                         std__mgr32__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane31_strm0_data        ;
  output                                        mgr32__std__lane31_strm0_data_valid  ;

  input                                         std__mgr32__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane31_strm1_data        ;
  output                                        mgr32__std__lane31_strm1_data_valid  ;

  input                                         std__mgr33__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane0_strm0_data        ;
  output                                        mgr33__std__lane0_strm0_data_valid  ;

  input                                         std__mgr33__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane0_strm1_data        ;
  output                                        mgr33__std__lane0_strm1_data_valid  ;

  input                                         std__mgr33__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane1_strm0_data        ;
  output                                        mgr33__std__lane1_strm0_data_valid  ;

  input                                         std__mgr33__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane1_strm1_data        ;
  output                                        mgr33__std__lane1_strm1_data_valid  ;

  input                                         std__mgr33__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane2_strm0_data        ;
  output                                        mgr33__std__lane2_strm0_data_valid  ;

  input                                         std__mgr33__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane2_strm1_data        ;
  output                                        mgr33__std__lane2_strm1_data_valid  ;

  input                                         std__mgr33__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane3_strm0_data        ;
  output                                        mgr33__std__lane3_strm0_data_valid  ;

  input                                         std__mgr33__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane3_strm1_data        ;
  output                                        mgr33__std__lane3_strm1_data_valid  ;

  input                                         std__mgr33__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane4_strm0_data        ;
  output                                        mgr33__std__lane4_strm0_data_valid  ;

  input                                         std__mgr33__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane4_strm1_data        ;
  output                                        mgr33__std__lane4_strm1_data_valid  ;

  input                                         std__mgr33__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane5_strm0_data        ;
  output                                        mgr33__std__lane5_strm0_data_valid  ;

  input                                         std__mgr33__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane5_strm1_data        ;
  output                                        mgr33__std__lane5_strm1_data_valid  ;

  input                                         std__mgr33__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane6_strm0_data        ;
  output                                        mgr33__std__lane6_strm0_data_valid  ;

  input                                         std__mgr33__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane6_strm1_data        ;
  output                                        mgr33__std__lane6_strm1_data_valid  ;

  input                                         std__mgr33__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane7_strm0_data        ;
  output                                        mgr33__std__lane7_strm0_data_valid  ;

  input                                         std__mgr33__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane7_strm1_data        ;
  output                                        mgr33__std__lane7_strm1_data_valid  ;

  input                                         std__mgr33__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane8_strm0_data        ;
  output                                        mgr33__std__lane8_strm0_data_valid  ;

  input                                         std__mgr33__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane8_strm1_data        ;
  output                                        mgr33__std__lane8_strm1_data_valid  ;

  input                                         std__mgr33__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane9_strm0_data        ;
  output                                        mgr33__std__lane9_strm0_data_valid  ;

  input                                         std__mgr33__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane9_strm1_data        ;
  output                                        mgr33__std__lane9_strm1_data_valid  ;

  input                                         std__mgr33__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane10_strm0_data        ;
  output                                        mgr33__std__lane10_strm0_data_valid  ;

  input                                         std__mgr33__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane10_strm1_data        ;
  output                                        mgr33__std__lane10_strm1_data_valid  ;

  input                                         std__mgr33__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane11_strm0_data        ;
  output                                        mgr33__std__lane11_strm0_data_valid  ;

  input                                         std__mgr33__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane11_strm1_data        ;
  output                                        mgr33__std__lane11_strm1_data_valid  ;

  input                                         std__mgr33__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane12_strm0_data        ;
  output                                        mgr33__std__lane12_strm0_data_valid  ;

  input                                         std__mgr33__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane12_strm1_data        ;
  output                                        mgr33__std__lane12_strm1_data_valid  ;

  input                                         std__mgr33__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane13_strm0_data        ;
  output                                        mgr33__std__lane13_strm0_data_valid  ;

  input                                         std__mgr33__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane13_strm1_data        ;
  output                                        mgr33__std__lane13_strm1_data_valid  ;

  input                                         std__mgr33__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane14_strm0_data        ;
  output                                        mgr33__std__lane14_strm0_data_valid  ;

  input                                         std__mgr33__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane14_strm1_data        ;
  output                                        mgr33__std__lane14_strm1_data_valid  ;

  input                                         std__mgr33__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane15_strm0_data        ;
  output                                        mgr33__std__lane15_strm0_data_valid  ;

  input                                         std__mgr33__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane15_strm1_data        ;
  output                                        mgr33__std__lane15_strm1_data_valid  ;

  input                                         std__mgr33__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane16_strm0_data        ;
  output                                        mgr33__std__lane16_strm0_data_valid  ;

  input                                         std__mgr33__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane16_strm1_data        ;
  output                                        mgr33__std__lane16_strm1_data_valid  ;

  input                                         std__mgr33__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane17_strm0_data        ;
  output                                        mgr33__std__lane17_strm0_data_valid  ;

  input                                         std__mgr33__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane17_strm1_data        ;
  output                                        mgr33__std__lane17_strm1_data_valid  ;

  input                                         std__mgr33__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane18_strm0_data        ;
  output                                        mgr33__std__lane18_strm0_data_valid  ;

  input                                         std__mgr33__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane18_strm1_data        ;
  output                                        mgr33__std__lane18_strm1_data_valid  ;

  input                                         std__mgr33__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane19_strm0_data        ;
  output                                        mgr33__std__lane19_strm0_data_valid  ;

  input                                         std__mgr33__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane19_strm1_data        ;
  output                                        mgr33__std__lane19_strm1_data_valid  ;

  input                                         std__mgr33__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane20_strm0_data        ;
  output                                        mgr33__std__lane20_strm0_data_valid  ;

  input                                         std__mgr33__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane20_strm1_data        ;
  output                                        mgr33__std__lane20_strm1_data_valid  ;

  input                                         std__mgr33__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane21_strm0_data        ;
  output                                        mgr33__std__lane21_strm0_data_valid  ;

  input                                         std__mgr33__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane21_strm1_data        ;
  output                                        mgr33__std__lane21_strm1_data_valid  ;

  input                                         std__mgr33__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane22_strm0_data        ;
  output                                        mgr33__std__lane22_strm0_data_valid  ;

  input                                         std__mgr33__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane22_strm1_data        ;
  output                                        mgr33__std__lane22_strm1_data_valid  ;

  input                                         std__mgr33__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane23_strm0_data        ;
  output                                        mgr33__std__lane23_strm0_data_valid  ;

  input                                         std__mgr33__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane23_strm1_data        ;
  output                                        mgr33__std__lane23_strm1_data_valid  ;

  input                                         std__mgr33__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane24_strm0_data        ;
  output                                        mgr33__std__lane24_strm0_data_valid  ;

  input                                         std__mgr33__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane24_strm1_data        ;
  output                                        mgr33__std__lane24_strm1_data_valid  ;

  input                                         std__mgr33__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane25_strm0_data        ;
  output                                        mgr33__std__lane25_strm0_data_valid  ;

  input                                         std__mgr33__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane25_strm1_data        ;
  output                                        mgr33__std__lane25_strm1_data_valid  ;

  input                                         std__mgr33__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane26_strm0_data        ;
  output                                        mgr33__std__lane26_strm0_data_valid  ;

  input                                         std__mgr33__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane26_strm1_data        ;
  output                                        mgr33__std__lane26_strm1_data_valid  ;

  input                                         std__mgr33__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane27_strm0_data        ;
  output                                        mgr33__std__lane27_strm0_data_valid  ;

  input                                         std__mgr33__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane27_strm1_data        ;
  output                                        mgr33__std__lane27_strm1_data_valid  ;

  input                                         std__mgr33__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane28_strm0_data        ;
  output                                        mgr33__std__lane28_strm0_data_valid  ;

  input                                         std__mgr33__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane28_strm1_data        ;
  output                                        mgr33__std__lane28_strm1_data_valid  ;

  input                                         std__mgr33__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane29_strm0_data        ;
  output                                        mgr33__std__lane29_strm0_data_valid  ;

  input                                         std__mgr33__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane29_strm1_data        ;
  output                                        mgr33__std__lane29_strm1_data_valid  ;

  input                                         std__mgr33__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane30_strm0_data        ;
  output                                        mgr33__std__lane30_strm0_data_valid  ;

  input                                         std__mgr33__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane30_strm1_data        ;
  output                                        mgr33__std__lane30_strm1_data_valid  ;

  input                                         std__mgr33__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane31_strm0_data        ;
  output                                        mgr33__std__lane31_strm0_data_valid  ;

  input                                         std__mgr33__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane31_strm1_data        ;
  output                                        mgr33__std__lane31_strm1_data_valid  ;

  input                                         std__mgr34__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane0_strm0_data        ;
  output                                        mgr34__std__lane0_strm0_data_valid  ;

  input                                         std__mgr34__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane0_strm1_data        ;
  output                                        mgr34__std__lane0_strm1_data_valid  ;

  input                                         std__mgr34__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane1_strm0_data        ;
  output                                        mgr34__std__lane1_strm0_data_valid  ;

  input                                         std__mgr34__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane1_strm1_data        ;
  output                                        mgr34__std__lane1_strm1_data_valid  ;

  input                                         std__mgr34__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane2_strm0_data        ;
  output                                        mgr34__std__lane2_strm0_data_valid  ;

  input                                         std__mgr34__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane2_strm1_data        ;
  output                                        mgr34__std__lane2_strm1_data_valid  ;

  input                                         std__mgr34__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane3_strm0_data        ;
  output                                        mgr34__std__lane3_strm0_data_valid  ;

  input                                         std__mgr34__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane3_strm1_data        ;
  output                                        mgr34__std__lane3_strm1_data_valid  ;

  input                                         std__mgr34__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane4_strm0_data        ;
  output                                        mgr34__std__lane4_strm0_data_valid  ;

  input                                         std__mgr34__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane4_strm1_data        ;
  output                                        mgr34__std__lane4_strm1_data_valid  ;

  input                                         std__mgr34__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane5_strm0_data        ;
  output                                        mgr34__std__lane5_strm0_data_valid  ;

  input                                         std__mgr34__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane5_strm1_data        ;
  output                                        mgr34__std__lane5_strm1_data_valid  ;

  input                                         std__mgr34__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane6_strm0_data        ;
  output                                        mgr34__std__lane6_strm0_data_valid  ;

  input                                         std__mgr34__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane6_strm1_data        ;
  output                                        mgr34__std__lane6_strm1_data_valid  ;

  input                                         std__mgr34__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane7_strm0_data        ;
  output                                        mgr34__std__lane7_strm0_data_valid  ;

  input                                         std__mgr34__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane7_strm1_data        ;
  output                                        mgr34__std__lane7_strm1_data_valid  ;

  input                                         std__mgr34__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane8_strm0_data        ;
  output                                        mgr34__std__lane8_strm0_data_valid  ;

  input                                         std__mgr34__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane8_strm1_data        ;
  output                                        mgr34__std__lane8_strm1_data_valid  ;

  input                                         std__mgr34__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane9_strm0_data        ;
  output                                        mgr34__std__lane9_strm0_data_valid  ;

  input                                         std__mgr34__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane9_strm1_data        ;
  output                                        mgr34__std__lane9_strm1_data_valid  ;

  input                                         std__mgr34__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane10_strm0_data        ;
  output                                        mgr34__std__lane10_strm0_data_valid  ;

  input                                         std__mgr34__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane10_strm1_data        ;
  output                                        mgr34__std__lane10_strm1_data_valid  ;

  input                                         std__mgr34__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane11_strm0_data        ;
  output                                        mgr34__std__lane11_strm0_data_valid  ;

  input                                         std__mgr34__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane11_strm1_data        ;
  output                                        mgr34__std__lane11_strm1_data_valid  ;

  input                                         std__mgr34__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane12_strm0_data        ;
  output                                        mgr34__std__lane12_strm0_data_valid  ;

  input                                         std__mgr34__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane12_strm1_data        ;
  output                                        mgr34__std__lane12_strm1_data_valid  ;

  input                                         std__mgr34__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane13_strm0_data        ;
  output                                        mgr34__std__lane13_strm0_data_valid  ;

  input                                         std__mgr34__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane13_strm1_data        ;
  output                                        mgr34__std__lane13_strm1_data_valid  ;

  input                                         std__mgr34__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane14_strm0_data        ;
  output                                        mgr34__std__lane14_strm0_data_valid  ;

  input                                         std__mgr34__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane14_strm1_data        ;
  output                                        mgr34__std__lane14_strm1_data_valid  ;

  input                                         std__mgr34__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane15_strm0_data        ;
  output                                        mgr34__std__lane15_strm0_data_valid  ;

  input                                         std__mgr34__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane15_strm1_data        ;
  output                                        mgr34__std__lane15_strm1_data_valid  ;

  input                                         std__mgr34__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane16_strm0_data        ;
  output                                        mgr34__std__lane16_strm0_data_valid  ;

  input                                         std__mgr34__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane16_strm1_data        ;
  output                                        mgr34__std__lane16_strm1_data_valid  ;

  input                                         std__mgr34__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane17_strm0_data        ;
  output                                        mgr34__std__lane17_strm0_data_valid  ;

  input                                         std__mgr34__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane17_strm1_data        ;
  output                                        mgr34__std__lane17_strm1_data_valid  ;

  input                                         std__mgr34__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane18_strm0_data        ;
  output                                        mgr34__std__lane18_strm0_data_valid  ;

  input                                         std__mgr34__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane18_strm1_data        ;
  output                                        mgr34__std__lane18_strm1_data_valid  ;

  input                                         std__mgr34__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane19_strm0_data        ;
  output                                        mgr34__std__lane19_strm0_data_valid  ;

  input                                         std__mgr34__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane19_strm1_data        ;
  output                                        mgr34__std__lane19_strm1_data_valid  ;

  input                                         std__mgr34__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane20_strm0_data        ;
  output                                        mgr34__std__lane20_strm0_data_valid  ;

  input                                         std__mgr34__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane20_strm1_data        ;
  output                                        mgr34__std__lane20_strm1_data_valid  ;

  input                                         std__mgr34__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane21_strm0_data        ;
  output                                        mgr34__std__lane21_strm0_data_valid  ;

  input                                         std__mgr34__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane21_strm1_data        ;
  output                                        mgr34__std__lane21_strm1_data_valid  ;

  input                                         std__mgr34__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane22_strm0_data        ;
  output                                        mgr34__std__lane22_strm0_data_valid  ;

  input                                         std__mgr34__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane22_strm1_data        ;
  output                                        mgr34__std__lane22_strm1_data_valid  ;

  input                                         std__mgr34__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane23_strm0_data        ;
  output                                        mgr34__std__lane23_strm0_data_valid  ;

  input                                         std__mgr34__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane23_strm1_data        ;
  output                                        mgr34__std__lane23_strm1_data_valid  ;

  input                                         std__mgr34__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane24_strm0_data        ;
  output                                        mgr34__std__lane24_strm0_data_valid  ;

  input                                         std__mgr34__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane24_strm1_data        ;
  output                                        mgr34__std__lane24_strm1_data_valid  ;

  input                                         std__mgr34__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane25_strm0_data        ;
  output                                        mgr34__std__lane25_strm0_data_valid  ;

  input                                         std__mgr34__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane25_strm1_data        ;
  output                                        mgr34__std__lane25_strm1_data_valid  ;

  input                                         std__mgr34__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane26_strm0_data        ;
  output                                        mgr34__std__lane26_strm0_data_valid  ;

  input                                         std__mgr34__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane26_strm1_data        ;
  output                                        mgr34__std__lane26_strm1_data_valid  ;

  input                                         std__mgr34__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane27_strm0_data        ;
  output                                        mgr34__std__lane27_strm0_data_valid  ;

  input                                         std__mgr34__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane27_strm1_data        ;
  output                                        mgr34__std__lane27_strm1_data_valid  ;

  input                                         std__mgr34__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane28_strm0_data        ;
  output                                        mgr34__std__lane28_strm0_data_valid  ;

  input                                         std__mgr34__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane28_strm1_data        ;
  output                                        mgr34__std__lane28_strm1_data_valid  ;

  input                                         std__mgr34__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane29_strm0_data        ;
  output                                        mgr34__std__lane29_strm0_data_valid  ;

  input                                         std__mgr34__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane29_strm1_data        ;
  output                                        mgr34__std__lane29_strm1_data_valid  ;

  input                                         std__mgr34__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane30_strm0_data        ;
  output                                        mgr34__std__lane30_strm0_data_valid  ;

  input                                         std__mgr34__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane30_strm1_data        ;
  output                                        mgr34__std__lane30_strm1_data_valid  ;

  input                                         std__mgr34__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane31_strm0_data        ;
  output                                        mgr34__std__lane31_strm0_data_valid  ;

  input                                         std__mgr34__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane31_strm1_data        ;
  output                                        mgr34__std__lane31_strm1_data_valid  ;

  input                                         std__mgr35__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane0_strm0_data        ;
  output                                        mgr35__std__lane0_strm0_data_valid  ;

  input                                         std__mgr35__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane0_strm1_data        ;
  output                                        mgr35__std__lane0_strm1_data_valid  ;

  input                                         std__mgr35__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane1_strm0_data        ;
  output                                        mgr35__std__lane1_strm0_data_valid  ;

  input                                         std__mgr35__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane1_strm1_data        ;
  output                                        mgr35__std__lane1_strm1_data_valid  ;

  input                                         std__mgr35__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane2_strm0_data        ;
  output                                        mgr35__std__lane2_strm0_data_valid  ;

  input                                         std__mgr35__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane2_strm1_data        ;
  output                                        mgr35__std__lane2_strm1_data_valid  ;

  input                                         std__mgr35__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane3_strm0_data        ;
  output                                        mgr35__std__lane3_strm0_data_valid  ;

  input                                         std__mgr35__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane3_strm1_data        ;
  output                                        mgr35__std__lane3_strm1_data_valid  ;

  input                                         std__mgr35__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane4_strm0_data        ;
  output                                        mgr35__std__lane4_strm0_data_valid  ;

  input                                         std__mgr35__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane4_strm1_data        ;
  output                                        mgr35__std__lane4_strm1_data_valid  ;

  input                                         std__mgr35__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane5_strm0_data        ;
  output                                        mgr35__std__lane5_strm0_data_valid  ;

  input                                         std__mgr35__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane5_strm1_data        ;
  output                                        mgr35__std__lane5_strm1_data_valid  ;

  input                                         std__mgr35__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane6_strm0_data        ;
  output                                        mgr35__std__lane6_strm0_data_valid  ;

  input                                         std__mgr35__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane6_strm1_data        ;
  output                                        mgr35__std__lane6_strm1_data_valid  ;

  input                                         std__mgr35__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane7_strm0_data        ;
  output                                        mgr35__std__lane7_strm0_data_valid  ;

  input                                         std__mgr35__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane7_strm1_data        ;
  output                                        mgr35__std__lane7_strm1_data_valid  ;

  input                                         std__mgr35__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane8_strm0_data        ;
  output                                        mgr35__std__lane8_strm0_data_valid  ;

  input                                         std__mgr35__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane8_strm1_data        ;
  output                                        mgr35__std__lane8_strm1_data_valid  ;

  input                                         std__mgr35__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane9_strm0_data        ;
  output                                        mgr35__std__lane9_strm0_data_valid  ;

  input                                         std__mgr35__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane9_strm1_data        ;
  output                                        mgr35__std__lane9_strm1_data_valid  ;

  input                                         std__mgr35__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane10_strm0_data        ;
  output                                        mgr35__std__lane10_strm0_data_valid  ;

  input                                         std__mgr35__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane10_strm1_data        ;
  output                                        mgr35__std__lane10_strm1_data_valid  ;

  input                                         std__mgr35__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane11_strm0_data        ;
  output                                        mgr35__std__lane11_strm0_data_valid  ;

  input                                         std__mgr35__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane11_strm1_data        ;
  output                                        mgr35__std__lane11_strm1_data_valid  ;

  input                                         std__mgr35__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane12_strm0_data        ;
  output                                        mgr35__std__lane12_strm0_data_valid  ;

  input                                         std__mgr35__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane12_strm1_data        ;
  output                                        mgr35__std__lane12_strm1_data_valid  ;

  input                                         std__mgr35__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane13_strm0_data        ;
  output                                        mgr35__std__lane13_strm0_data_valid  ;

  input                                         std__mgr35__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane13_strm1_data        ;
  output                                        mgr35__std__lane13_strm1_data_valid  ;

  input                                         std__mgr35__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane14_strm0_data        ;
  output                                        mgr35__std__lane14_strm0_data_valid  ;

  input                                         std__mgr35__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane14_strm1_data        ;
  output                                        mgr35__std__lane14_strm1_data_valid  ;

  input                                         std__mgr35__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane15_strm0_data        ;
  output                                        mgr35__std__lane15_strm0_data_valid  ;

  input                                         std__mgr35__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane15_strm1_data        ;
  output                                        mgr35__std__lane15_strm1_data_valid  ;

  input                                         std__mgr35__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane16_strm0_data        ;
  output                                        mgr35__std__lane16_strm0_data_valid  ;

  input                                         std__mgr35__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane16_strm1_data        ;
  output                                        mgr35__std__lane16_strm1_data_valid  ;

  input                                         std__mgr35__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane17_strm0_data        ;
  output                                        mgr35__std__lane17_strm0_data_valid  ;

  input                                         std__mgr35__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane17_strm1_data        ;
  output                                        mgr35__std__lane17_strm1_data_valid  ;

  input                                         std__mgr35__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane18_strm0_data        ;
  output                                        mgr35__std__lane18_strm0_data_valid  ;

  input                                         std__mgr35__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane18_strm1_data        ;
  output                                        mgr35__std__lane18_strm1_data_valid  ;

  input                                         std__mgr35__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane19_strm0_data        ;
  output                                        mgr35__std__lane19_strm0_data_valid  ;

  input                                         std__mgr35__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane19_strm1_data        ;
  output                                        mgr35__std__lane19_strm1_data_valid  ;

  input                                         std__mgr35__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane20_strm0_data        ;
  output                                        mgr35__std__lane20_strm0_data_valid  ;

  input                                         std__mgr35__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane20_strm1_data        ;
  output                                        mgr35__std__lane20_strm1_data_valid  ;

  input                                         std__mgr35__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane21_strm0_data        ;
  output                                        mgr35__std__lane21_strm0_data_valid  ;

  input                                         std__mgr35__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane21_strm1_data        ;
  output                                        mgr35__std__lane21_strm1_data_valid  ;

  input                                         std__mgr35__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane22_strm0_data        ;
  output                                        mgr35__std__lane22_strm0_data_valid  ;

  input                                         std__mgr35__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane22_strm1_data        ;
  output                                        mgr35__std__lane22_strm1_data_valid  ;

  input                                         std__mgr35__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane23_strm0_data        ;
  output                                        mgr35__std__lane23_strm0_data_valid  ;

  input                                         std__mgr35__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane23_strm1_data        ;
  output                                        mgr35__std__lane23_strm1_data_valid  ;

  input                                         std__mgr35__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane24_strm0_data        ;
  output                                        mgr35__std__lane24_strm0_data_valid  ;

  input                                         std__mgr35__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane24_strm1_data        ;
  output                                        mgr35__std__lane24_strm1_data_valid  ;

  input                                         std__mgr35__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane25_strm0_data        ;
  output                                        mgr35__std__lane25_strm0_data_valid  ;

  input                                         std__mgr35__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane25_strm1_data        ;
  output                                        mgr35__std__lane25_strm1_data_valid  ;

  input                                         std__mgr35__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane26_strm0_data        ;
  output                                        mgr35__std__lane26_strm0_data_valid  ;

  input                                         std__mgr35__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane26_strm1_data        ;
  output                                        mgr35__std__lane26_strm1_data_valid  ;

  input                                         std__mgr35__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane27_strm0_data        ;
  output                                        mgr35__std__lane27_strm0_data_valid  ;

  input                                         std__mgr35__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane27_strm1_data        ;
  output                                        mgr35__std__lane27_strm1_data_valid  ;

  input                                         std__mgr35__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane28_strm0_data        ;
  output                                        mgr35__std__lane28_strm0_data_valid  ;

  input                                         std__mgr35__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane28_strm1_data        ;
  output                                        mgr35__std__lane28_strm1_data_valid  ;

  input                                         std__mgr35__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane29_strm0_data        ;
  output                                        mgr35__std__lane29_strm0_data_valid  ;

  input                                         std__mgr35__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane29_strm1_data        ;
  output                                        mgr35__std__lane29_strm1_data_valid  ;

  input                                         std__mgr35__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane30_strm0_data        ;
  output                                        mgr35__std__lane30_strm0_data_valid  ;

  input                                         std__mgr35__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane30_strm1_data        ;
  output                                        mgr35__std__lane30_strm1_data_valid  ;

  input                                         std__mgr35__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane31_strm0_data        ;
  output                                        mgr35__std__lane31_strm0_data_valid  ;

  input                                         std__mgr35__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane31_strm1_data        ;
  output                                        mgr35__std__lane31_strm1_data_valid  ;

  input                                         std__mgr36__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane0_strm0_data        ;
  output                                        mgr36__std__lane0_strm0_data_valid  ;

  input                                         std__mgr36__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane0_strm1_data        ;
  output                                        mgr36__std__lane0_strm1_data_valid  ;

  input                                         std__mgr36__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane1_strm0_data        ;
  output                                        mgr36__std__lane1_strm0_data_valid  ;

  input                                         std__mgr36__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane1_strm1_data        ;
  output                                        mgr36__std__lane1_strm1_data_valid  ;

  input                                         std__mgr36__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane2_strm0_data        ;
  output                                        mgr36__std__lane2_strm0_data_valid  ;

  input                                         std__mgr36__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane2_strm1_data        ;
  output                                        mgr36__std__lane2_strm1_data_valid  ;

  input                                         std__mgr36__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane3_strm0_data        ;
  output                                        mgr36__std__lane3_strm0_data_valid  ;

  input                                         std__mgr36__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane3_strm1_data        ;
  output                                        mgr36__std__lane3_strm1_data_valid  ;

  input                                         std__mgr36__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane4_strm0_data        ;
  output                                        mgr36__std__lane4_strm0_data_valid  ;

  input                                         std__mgr36__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane4_strm1_data        ;
  output                                        mgr36__std__lane4_strm1_data_valid  ;

  input                                         std__mgr36__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane5_strm0_data        ;
  output                                        mgr36__std__lane5_strm0_data_valid  ;

  input                                         std__mgr36__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane5_strm1_data        ;
  output                                        mgr36__std__lane5_strm1_data_valid  ;

  input                                         std__mgr36__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane6_strm0_data        ;
  output                                        mgr36__std__lane6_strm0_data_valid  ;

  input                                         std__mgr36__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane6_strm1_data        ;
  output                                        mgr36__std__lane6_strm1_data_valid  ;

  input                                         std__mgr36__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane7_strm0_data        ;
  output                                        mgr36__std__lane7_strm0_data_valid  ;

  input                                         std__mgr36__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane7_strm1_data        ;
  output                                        mgr36__std__lane7_strm1_data_valid  ;

  input                                         std__mgr36__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane8_strm0_data        ;
  output                                        mgr36__std__lane8_strm0_data_valid  ;

  input                                         std__mgr36__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane8_strm1_data        ;
  output                                        mgr36__std__lane8_strm1_data_valid  ;

  input                                         std__mgr36__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane9_strm0_data        ;
  output                                        mgr36__std__lane9_strm0_data_valid  ;

  input                                         std__mgr36__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane9_strm1_data        ;
  output                                        mgr36__std__lane9_strm1_data_valid  ;

  input                                         std__mgr36__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane10_strm0_data        ;
  output                                        mgr36__std__lane10_strm0_data_valid  ;

  input                                         std__mgr36__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane10_strm1_data        ;
  output                                        mgr36__std__lane10_strm1_data_valid  ;

  input                                         std__mgr36__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane11_strm0_data        ;
  output                                        mgr36__std__lane11_strm0_data_valid  ;

  input                                         std__mgr36__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane11_strm1_data        ;
  output                                        mgr36__std__lane11_strm1_data_valid  ;

  input                                         std__mgr36__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane12_strm0_data        ;
  output                                        mgr36__std__lane12_strm0_data_valid  ;

  input                                         std__mgr36__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane12_strm1_data        ;
  output                                        mgr36__std__lane12_strm1_data_valid  ;

  input                                         std__mgr36__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane13_strm0_data        ;
  output                                        mgr36__std__lane13_strm0_data_valid  ;

  input                                         std__mgr36__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane13_strm1_data        ;
  output                                        mgr36__std__lane13_strm1_data_valid  ;

  input                                         std__mgr36__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane14_strm0_data        ;
  output                                        mgr36__std__lane14_strm0_data_valid  ;

  input                                         std__mgr36__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane14_strm1_data        ;
  output                                        mgr36__std__lane14_strm1_data_valid  ;

  input                                         std__mgr36__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane15_strm0_data        ;
  output                                        mgr36__std__lane15_strm0_data_valid  ;

  input                                         std__mgr36__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane15_strm1_data        ;
  output                                        mgr36__std__lane15_strm1_data_valid  ;

  input                                         std__mgr36__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane16_strm0_data        ;
  output                                        mgr36__std__lane16_strm0_data_valid  ;

  input                                         std__mgr36__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane16_strm1_data        ;
  output                                        mgr36__std__lane16_strm1_data_valid  ;

  input                                         std__mgr36__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane17_strm0_data        ;
  output                                        mgr36__std__lane17_strm0_data_valid  ;

  input                                         std__mgr36__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane17_strm1_data        ;
  output                                        mgr36__std__lane17_strm1_data_valid  ;

  input                                         std__mgr36__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane18_strm0_data        ;
  output                                        mgr36__std__lane18_strm0_data_valid  ;

  input                                         std__mgr36__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane18_strm1_data        ;
  output                                        mgr36__std__lane18_strm1_data_valid  ;

  input                                         std__mgr36__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane19_strm0_data        ;
  output                                        mgr36__std__lane19_strm0_data_valid  ;

  input                                         std__mgr36__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane19_strm1_data        ;
  output                                        mgr36__std__lane19_strm1_data_valid  ;

  input                                         std__mgr36__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane20_strm0_data        ;
  output                                        mgr36__std__lane20_strm0_data_valid  ;

  input                                         std__mgr36__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane20_strm1_data        ;
  output                                        mgr36__std__lane20_strm1_data_valid  ;

  input                                         std__mgr36__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane21_strm0_data        ;
  output                                        mgr36__std__lane21_strm0_data_valid  ;

  input                                         std__mgr36__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane21_strm1_data        ;
  output                                        mgr36__std__lane21_strm1_data_valid  ;

  input                                         std__mgr36__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane22_strm0_data        ;
  output                                        mgr36__std__lane22_strm0_data_valid  ;

  input                                         std__mgr36__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane22_strm1_data        ;
  output                                        mgr36__std__lane22_strm1_data_valid  ;

  input                                         std__mgr36__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane23_strm0_data        ;
  output                                        mgr36__std__lane23_strm0_data_valid  ;

  input                                         std__mgr36__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane23_strm1_data        ;
  output                                        mgr36__std__lane23_strm1_data_valid  ;

  input                                         std__mgr36__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane24_strm0_data        ;
  output                                        mgr36__std__lane24_strm0_data_valid  ;

  input                                         std__mgr36__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane24_strm1_data        ;
  output                                        mgr36__std__lane24_strm1_data_valid  ;

  input                                         std__mgr36__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane25_strm0_data        ;
  output                                        mgr36__std__lane25_strm0_data_valid  ;

  input                                         std__mgr36__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane25_strm1_data        ;
  output                                        mgr36__std__lane25_strm1_data_valid  ;

  input                                         std__mgr36__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane26_strm0_data        ;
  output                                        mgr36__std__lane26_strm0_data_valid  ;

  input                                         std__mgr36__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane26_strm1_data        ;
  output                                        mgr36__std__lane26_strm1_data_valid  ;

  input                                         std__mgr36__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane27_strm0_data        ;
  output                                        mgr36__std__lane27_strm0_data_valid  ;

  input                                         std__mgr36__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane27_strm1_data        ;
  output                                        mgr36__std__lane27_strm1_data_valid  ;

  input                                         std__mgr36__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane28_strm0_data        ;
  output                                        mgr36__std__lane28_strm0_data_valid  ;

  input                                         std__mgr36__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane28_strm1_data        ;
  output                                        mgr36__std__lane28_strm1_data_valid  ;

  input                                         std__mgr36__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane29_strm0_data        ;
  output                                        mgr36__std__lane29_strm0_data_valid  ;

  input                                         std__mgr36__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane29_strm1_data        ;
  output                                        mgr36__std__lane29_strm1_data_valid  ;

  input                                         std__mgr36__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane30_strm0_data        ;
  output                                        mgr36__std__lane30_strm0_data_valid  ;

  input                                         std__mgr36__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane30_strm1_data        ;
  output                                        mgr36__std__lane30_strm1_data_valid  ;

  input                                         std__mgr36__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane31_strm0_data        ;
  output                                        mgr36__std__lane31_strm0_data_valid  ;

  input                                         std__mgr36__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane31_strm1_data        ;
  output                                        mgr36__std__lane31_strm1_data_valid  ;

  input                                         std__mgr37__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane0_strm0_data        ;
  output                                        mgr37__std__lane0_strm0_data_valid  ;

  input                                         std__mgr37__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane0_strm1_data        ;
  output                                        mgr37__std__lane0_strm1_data_valid  ;

  input                                         std__mgr37__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane1_strm0_data        ;
  output                                        mgr37__std__lane1_strm0_data_valid  ;

  input                                         std__mgr37__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane1_strm1_data        ;
  output                                        mgr37__std__lane1_strm1_data_valid  ;

  input                                         std__mgr37__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane2_strm0_data        ;
  output                                        mgr37__std__lane2_strm0_data_valid  ;

  input                                         std__mgr37__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane2_strm1_data        ;
  output                                        mgr37__std__lane2_strm1_data_valid  ;

  input                                         std__mgr37__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane3_strm0_data        ;
  output                                        mgr37__std__lane3_strm0_data_valid  ;

  input                                         std__mgr37__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane3_strm1_data        ;
  output                                        mgr37__std__lane3_strm1_data_valid  ;

  input                                         std__mgr37__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane4_strm0_data        ;
  output                                        mgr37__std__lane4_strm0_data_valid  ;

  input                                         std__mgr37__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane4_strm1_data        ;
  output                                        mgr37__std__lane4_strm1_data_valid  ;

  input                                         std__mgr37__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane5_strm0_data        ;
  output                                        mgr37__std__lane5_strm0_data_valid  ;

  input                                         std__mgr37__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane5_strm1_data        ;
  output                                        mgr37__std__lane5_strm1_data_valid  ;

  input                                         std__mgr37__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane6_strm0_data        ;
  output                                        mgr37__std__lane6_strm0_data_valid  ;

  input                                         std__mgr37__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane6_strm1_data        ;
  output                                        mgr37__std__lane6_strm1_data_valid  ;

  input                                         std__mgr37__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane7_strm0_data        ;
  output                                        mgr37__std__lane7_strm0_data_valid  ;

  input                                         std__mgr37__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane7_strm1_data        ;
  output                                        mgr37__std__lane7_strm1_data_valid  ;

  input                                         std__mgr37__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane8_strm0_data        ;
  output                                        mgr37__std__lane8_strm0_data_valid  ;

  input                                         std__mgr37__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane8_strm1_data        ;
  output                                        mgr37__std__lane8_strm1_data_valid  ;

  input                                         std__mgr37__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane9_strm0_data        ;
  output                                        mgr37__std__lane9_strm0_data_valid  ;

  input                                         std__mgr37__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane9_strm1_data        ;
  output                                        mgr37__std__lane9_strm1_data_valid  ;

  input                                         std__mgr37__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane10_strm0_data        ;
  output                                        mgr37__std__lane10_strm0_data_valid  ;

  input                                         std__mgr37__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane10_strm1_data        ;
  output                                        mgr37__std__lane10_strm1_data_valid  ;

  input                                         std__mgr37__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane11_strm0_data        ;
  output                                        mgr37__std__lane11_strm0_data_valid  ;

  input                                         std__mgr37__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane11_strm1_data        ;
  output                                        mgr37__std__lane11_strm1_data_valid  ;

  input                                         std__mgr37__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane12_strm0_data        ;
  output                                        mgr37__std__lane12_strm0_data_valid  ;

  input                                         std__mgr37__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane12_strm1_data        ;
  output                                        mgr37__std__lane12_strm1_data_valid  ;

  input                                         std__mgr37__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane13_strm0_data        ;
  output                                        mgr37__std__lane13_strm0_data_valid  ;

  input                                         std__mgr37__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane13_strm1_data        ;
  output                                        mgr37__std__lane13_strm1_data_valid  ;

  input                                         std__mgr37__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane14_strm0_data        ;
  output                                        mgr37__std__lane14_strm0_data_valid  ;

  input                                         std__mgr37__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane14_strm1_data        ;
  output                                        mgr37__std__lane14_strm1_data_valid  ;

  input                                         std__mgr37__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane15_strm0_data        ;
  output                                        mgr37__std__lane15_strm0_data_valid  ;

  input                                         std__mgr37__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane15_strm1_data        ;
  output                                        mgr37__std__lane15_strm1_data_valid  ;

  input                                         std__mgr37__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane16_strm0_data        ;
  output                                        mgr37__std__lane16_strm0_data_valid  ;

  input                                         std__mgr37__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane16_strm1_data        ;
  output                                        mgr37__std__lane16_strm1_data_valid  ;

  input                                         std__mgr37__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane17_strm0_data        ;
  output                                        mgr37__std__lane17_strm0_data_valid  ;

  input                                         std__mgr37__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane17_strm1_data        ;
  output                                        mgr37__std__lane17_strm1_data_valid  ;

  input                                         std__mgr37__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane18_strm0_data        ;
  output                                        mgr37__std__lane18_strm0_data_valid  ;

  input                                         std__mgr37__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane18_strm1_data        ;
  output                                        mgr37__std__lane18_strm1_data_valid  ;

  input                                         std__mgr37__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane19_strm0_data        ;
  output                                        mgr37__std__lane19_strm0_data_valid  ;

  input                                         std__mgr37__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane19_strm1_data        ;
  output                                        mgr37__std__lane19_strm1_data_valid  ;

  input                                         std__mgr37__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane20_strm0_data        ;
  output                                        mgr37__std__lane20_strm0_data_valid  ;

  input                                         std__mgr37__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane20_strm1_data        ;
  output                                        mgr37__std__lane20_strm1_data_valid  ;

  input                                         std__mgr37__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane21_strm0_data        ;
  output                                        mgr37__std__lane21_strm0_data_valid  ;

  input                                         std__mgr37__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane21_strm1_data        ;
  output                                        mgr37__std__lane21_strm1_data_valid  ;

  input                                         std__mgr37__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane22_strm0_data        ;
  output                                        mgr37__std__lane22_strm0_data_valid  ;

  input                                         std__mgr37__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane22_strm1_data        ;
  output                                        mgr37__std__lane22_strm1_data_valid  ;

  input                                         std__mgr37__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane23_strm0_data        ;
  output                                        mgr37__std__lane23_strm0_data_valid  ;

  input                                         std__mgr37__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane23_strm1_data        ;
  output                                        mgr37__std__lane23_strm1_data_valid  ;

  input                                         std__mgr37__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane24_strm0_data        ;
  output                                        mgr37__std__lane24_strm0_data_valid  ;

  input                                         std__mgr37__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane24_strm1_data        ;
  output                                        mgr37__std__lane24_strm1_data_valid  ;

  input                                         std__mgr37__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane25_strm0_data        ;
  output                                        mgr37__std__lane25_strm0_data_valid  ;

  input                                         std__mgr37__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane25_strm1_data        ;
  output                                        mgr37__std__lane25_strm1_data_valid  ;

  input                                         std__mgr37__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane26_strm0_data        ;
  output                                        mgr37__std__lane26_strm0_data_valid  ;

  input                                         std__mgr37__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane26_strm1_data        ;
  output                                        mgr37__std__lane26_strm1_data_valid  ;

  input                                         std__mgr37__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane27_strm0_data        ;
  output                                        mgr37__std__lane27_strm0_data_valid  ;

  input                                         std__mgr37__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane27_strm1_data        ;
  output                                        mgr37__std__lane27_strm1_data_valid  ;

  input                                         std__mgr37__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane28_strm0_data        ;
  output                                        mgr37__std__lane28_strm0_data_valid  ;

  input                                         std__mgr37__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane28_strm1_data        ;
  output                                        mgr37__std__lane28_strm1_data_valid  ;

  input                                         std__mgr37__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane29_strm0_data        ;
  output                                        mgr37__std__lane29_strm0_data_valid  ;

  input                                         std__mgr37__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane29_strm1_data        ;
  output                                        mgr37__std__lane29_strm1_data_valid  ;

  input                                         std__mgr37__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane30_strm0_data        ;
  output                                        mgr37__std__lane30_strm0_data_valid  ;

  input                                         std__mgr37__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane30_strm1_data        ;
  output                                        mgr37__std__lane30_strm1_data_valid  ;

  input                                         std__mgr37__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane31_strm0_data        ;
  output                                        mgr37__std__lane31_strm0_data_valid  ;

  input                                         std__mgr37__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane31_strm1_data        ;
  output                                        mgr37__std__lane31_strm1_data_valid  ;

  input                                         std__mgr38__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane0_strm0_data        ;
  output                                        mgr38__std__lane0_strm0_data_valid  ;

  input                                         std__mgr38__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane0_strm1_data        ;
  output                                        mgr38__std__lane0_strm1_data_valid  ;

  input                                         std__mgr38__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane1_strm0_data        ;
  output                                        mgr38__std__lane1_strm0_data_valid  ;

  input                                         std__mgr38__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane1_strm1_data        ;
  output                                        mgr38__std__lane1_strm1_data_valid  ;

  input                                         std__mgr38__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane2_strm0_data        ;
  output                                        mgr38__std__lane2_strm0_data_valid  ;

  input                                         std__mgr38__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane2_strm1_data        ;
  output                                        mgr38__std__lane2_strm1_data_valid  ;

  input                                         std__mgr38__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane3_strm0_data        ;
  output                                        mgr38__std__lane3_strm0_data_valid  ;

  input                                         std__mgr38__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane3_strm1_data        ;
  output                                        mgr38__std__lane3_strm1_data_valid  ;

  input                                         std__mgr38__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane4_strm0_data        ;
  output                                        mgr38__std__lane4_strm0_data_valid  ;

  input                                         std__mgr38__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane4_strm1_data        ;
  output                                        mgr38__std__lane4_strm1_data_valid  ;

  input                                         std__mgr38__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane5_strm0_data        ;
  output                                        mgr38__std__lane5_strm0_data_valid  ;

  input                                         std__mgr38__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane5_strm1_data        ;
  output                                        mgr38__std__lane5_strm1_data_valid  ;

  input                                         std__mgr38__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane6_strm0_data        ;
  output                                        mgr38__std__lane6_strm0_data_valid  ;

  input                                         std__mgr38__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane6_strm1_data        ;
  output                                        mgr38__std__lane6_strm1_data_valid  ;

  input                                         std__mgr38__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane7_strm0_data        ;
  output                                        mgr38__std__lane7_strm0_data_valid  ;

  input                                         std__mgr38__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane7_strm1_data        ;
  output                                        mgr38__std__lane7_strm1_data_valid  ;

  input                                         std__mgr38__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane8_strm0_data        ;
  output                                        mgr38__std__lane8_strm0_data_valid  ;

  input                                         std__mgr38__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane8_strm1_data        ;
  output                                        mgr38__std__lane8_strm1_data_valid  ;

  input                                         std__mgr38__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane9_strm0_data        ;
  output                                        mgr38__std__lane9_strm0_data_valid  ;

  input                                         std__mgr38__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane9_strm1_data        ;
  output                                        mgr38__std__lane9_strm1_data_valid  ;

  input                                         std__mgr38__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane10_strm0_data        ;
  output                                        mgr38__std__lane10_strm0_data_valid  ;

  input                                         std__mgr38__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane10_strm1_data        ;
  output                                        mgr38__std__lane10_strm1_data_valid  ;

  input                                         std__mgr38__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane11_strm0_data        ;
  output                                        mgr38__std__lane11_strm0_data_valid  ;

  input                                         std__mgr38__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane11_strm1_data        ;
  output                                        mgr38__std__lane11_strm1_data_valid  ;

  input                                         std__mgr38__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane12_strm0_data        ;
  output                                        mgr38__std__lane12_strm0_data_valid  ;

  input                                         std__mgr38__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane12_strm1_data        ;
  output                                        mgr38__std__lane12_strm1_data_valid  ;

  input                                         std__mgr38__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane13_strm0_data        ;
  output                                        mgr38__std__lane13_strm0_data_valid  ;

  input                                         std__mgr38__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane13_strm1_data        ;
  output                                        mgr38__std__lane13_strm1_data_valid  ;

  input                                         std__mgr38__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane14_strm0_data        ;
  output                                        mgr38__std__lane14_strm0_data_valid  ;

  input                                         std__mgr38__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane14_strm1_data        ;
  output                                        mgr38__std__lane14_strm1_data_valid  ;

  input                                         std__mgr38__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane15_strm0_data        ;
  output                                        mgr38__std__lane15_strm0_data_valid  ;

  input                                         std__mgr38__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane15_strm1_data        ;
  output                                        mgr38__std__lane15_strm1_data_valid  ;

  input                                         std__mgr38__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane16_strm0_data        ;
  output                                        mgr38__std__lane16_strm0_data_valid  ;

  input                                         std__mgr38__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane16_strm1_data        ;
  output                                        mgr38__std__lane16_strm1_data_valid  ;

  input                                         std__mgr38__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane17_strm0_data        ;
  output                                        mgr38__std__lane17_strm0_data_valid  ;

  input                                         std__mgr38__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane17_strm1_data        ;
  output                                        mgr38__std__lane17_strm1_data_valid  ;

  input                                         std__mgr38__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane18_strm0_data        ;
  output                                        mgr38__std__lane18_strm0_data_valid  ;

  input                                         std__mgr38__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane18_strm1_data        ;
  output                                        mgr38__std__lane18_strm1_data_valid  ;

  input                                         std__mgr38__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane19_strm0_data        ;
  output                                        mgr38__std__lane19_strm0_data_valid  ;

  input                                         std__mgr38__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane19_strm1_data        ;
  output                                        mgr38__std__lane19_strm1_data_valid  ;

  input                                         std__mgr38__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane20_strm0_data        ;
  output                                        mgr38__std__lane20_strm0_data_valid  ;

  input                                         std__mgr38__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane20_strm1_data        ;
  output                                        mgr38__std__lane20_strm1_data_valid  ;

  input                                         std__mgr38__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane21_strm0_data        ;
  output                                        mgr38__std__lane21_strm0_data_valid  ;

  input                                         std__mgr38__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane21_strm1_data        ;
  output                                        mgr38__std__lane21_strm1_data_valid  ;

  input                                         std__mgr38__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane22_strm0_data        ;
  output                                        mgr38__std__lane22_strm0_data_valid  ;

  input                                         std__mgr38__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane22_strm1_data        ;
  output                                        mgr38__std__lane22_strm1_data_valid  ;

  input                                         std__mgr38__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane23_strm0_data        ;
  output                                        mgr38__std__lane23_strm0_data_valid  ;

  input                                         std__mgr38__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane23_strm1_data        ;
  output                                        mgr38__std__lane23_strm1_data_valid  ;

  input                                         std__mgr38__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane24_strm0_data        ;
  output                                        mgr38__std__lane24_strm0_data_valid  ;

  input                                         std__mgr38__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane24_strm1_data        ;
  output                                        mgr38__std__lane24_strm1_data_valid  ;

  input                                         std__mgr38__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane25_strm0_data        ;
  output                                        mgr38__std__lane25_strm0_data_valid  ;

  input                                         std__mgr38__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane25_strm1_data        ;
  output                                        mgr38__std__lane25_strm1_data_valid  ;

  input                                         std__mgr38__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane26_strm0_data        ;
  output                                        mgr38__std__lane26_strm0_data_valid  ;

  input                                         std__mgr38__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane26_strm1_data        ;
  output                                        mgr38__std__lane26_strm1_data_valid  ;

  input                                         std__mgr38__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane27_strm0_data        ;
  output                                        mgr38__std__lane27_strm0_data_valid  ;

  input                                         std__mgr38__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane27_strm1_data        ;
  output                                        mgr38__std__lane27_strm1_data_valid  ;

  input                                         std__mgr38__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane28_strm0_data        ;
  output                                        mgr38__std__lane28_strm0_data_valid  ;

  input                                         std__mgr38__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane28_strm1_data        ;
  output                                        mgr38__std__lane28_strm1_data_valid  ;

  input                                         std__mgr38__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane29_strm0_data        ;
  output                                        mgr38__std__lane29_strm0_data_valid  ;

  input                                         std__mgr38__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane29_strm1_data        ;
  output                                        mgr38__std__lane29_strm1_data_valid  ;

  input                                         std__mgr38__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane30_strm0_data        ;
  output                                        mgr38__std__lane30_strm0_data_valid  ;

  input                                         std__mgr38__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane30_strm1_data        ;
  output                                        mgr38__std__lane30_strm1_data_valid  ;

  input                                         std__mgr38__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane31_strm0_data        ;
  output                                        mgr38__std__lane31_strm0_data_valid  ;

  input                                         std__mgr38__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane31_strm1_data        ;
  output                                        mgr38__std__lane31_strm1_data_valid  ;

  input                                         std__mgr39__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane0_strm0_data        ;
  output                                        mgr39__std__lane0_strm0_data_valid  ;

  input                                         std__mgr39__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane0_strm1_data        ;
  output                                        mgr39__std__lane0_strm1_data_valid  ;

  input                                         std__mgr39__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane1_strm0_data        ;
  output                                        mgr39__std__lane1_strm0_data_valid  ;

  input                                         std__mgr39__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane1_strm1_data        ;
  output                                        mgr39__std__lane1_strm1_data_valid  ;

  input                                         std__mgr39__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane2_strm0_data        ;
  output                                        mgr39__std__lane2_strm0_data_valid  ;

  input                                         std__mgr39__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane2_strm1_data        ;
  output                                        mgr39__std__lane2_strm1_data_valid  ;

  input                                         std__mgr39__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane3_strm0_data        ;
  output                                        mgr39__std__lane3_strm0_data_valid  ;

  input                                         std__mgr39__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane3_strm1_data        ;
  output                                        mgr39__std__lane3_strm1_data_valid  ;

  input                                         std__mgr39__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane4_strm0_data        ;
  output                                        mgr39__std__lane4_strm0_data_valid  ;

  input                                         std__mgr39__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane4_strm1_data        ;
  output                                        mgr39__std__lane4_strm1_data_valid  ;

  input                                         std__mgr39__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane5_strm0_data        ;
  output                                        mgr39__std__lane5_strm0_data_valid  ;

  input                                         std__mgr39__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane5_strm1_data        ;
  output                                        mgr39__std__lane5_strm1_data_valid  ;

  input                                         std__mgr39__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane6_strm0_data        ;
  output                                        mgr39__std__lane6_strm0_data_valid  ;

  input                                         std__mgr39__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane6_strm1_data        ;
  output                                        mgr39__std__lane6_strm1_data_valid  ;

  input                                         std__mgr39__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane7_strm0_data        ;
  output                                        mgr39__std__lane7_strm0_data_valid  ;

  input                                         std__mgr39__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane7_strm1_data        ;
  output                                        mgr39__std__lane7_strm1_data_valid  ;

  input                                         std__mgr39__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane8_strm0_data        ;
  output                                        mgr39__std__lane8_strm0_data_valid  ;

  input                                         std__mgr39__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane8_strm1_data        ;
  output                                        mgr39__std__lane8_strm1_data_valid  ;

  input                                         std__mgr39__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane9_strm0_data        ;
  output                                        mgr39__std__lane9_strm0_data_valid  ;

  input                                         std__mgr39__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane9_strm1_data        ;
  output                                        mgr39__std__lane9_strm1_data_valid  ;

  input                                         std__mgr39__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane10_strm0_data        ;
  output                                        mgr39__std__lane10_strm0_data_valid  ;

  input                                         std__mgr39__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane10_strm1_data        ;
  output                                        mgr39__std__lane10_strm1_data_valid  ;

  input                                         std__mgr39__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane11_strm0_data        ;
  output                                        mgr39__std__lane11_strm0_data_valid  ;

  input                                         std__mgr39__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane11_strm1_data        ;
  output                                        mgr39__std__lane11_strm1_data_valid  ;

  input                                         std__mgr39__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane12_strm0_data        ;
  output                                        mgr39__std__lane12_strm0_data_valid  ;

  input                                         std__mgr39__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane12_strm1_data        ;
  output                                        mgr39__std__lane12_strm1_data_valid  ;

  input                                         std__mgr39__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane13_strm0_data        ;
  output                                        mgr39__std__lane13_strm0_data_valid  ;

  input                                         std__mgr39__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane13_strm1_data        ;
  output                                        mgr39__std__lane13_strm1_data_valid  ;

  input                                         std__mgr39__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane14_strm0_data        ;
  output                                        mgr39__std__lane14_strm0_data_valid  ;

  input                                         std__mgr39__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane14_strm1_data        ;
  output                                        mgr39__std__lane14_strm1_data_valid  ;

  input                                         std__mgr39__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane15_strm0_data        ;
  output                                        mgr39__std__lane15_strm0_data_valid  ;

  input                                         std__mgr39__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane15_strm1_data        ;
  output                                        mgr39__std__lane15_strm1_data_valid  ;

  input                                         std__mgr39__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane16_strm0_data        ;
  output                                        mgr39__std__lane16_strm0_data_valid  ;

  input                                         std__mgr39__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane16_strm1_data        ;
  output                                        mgr39__std__lane16_strm1_data_valid  ;

  input                                         std__mgr39__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane17_strm0_data        ;
  output                                        mgr39__std__lane17_strm0_data_valid  ;

  input                                         std__mgr39__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane17_strm1_data        ;
  output                                        mgr39__std__lane17_strm1_data_valid  ;

  input                                         std__mgr39__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane18_strm0_data        ;
  output                                        mgr39__std__lane18_strm0_data_valid  ;

  input                                         std__mgr39__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane18_strm1_data        ;
  output                                        mgr39__std__lane18_strm1_data_valid  ;

  input                                         std__mgr39__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane19_strm0_data        ;
  output                                        mgr39__std__lane19_strm0_data_valid  ;

  input                                         std__mgr39__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane19_strm1_data        ;
  output                                        mgr39__std__lane19_strm1_data_valid  ;

  input                                         std__mgr39__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane20_strm0_data        ;
  output                                        mgr39__std__lane20_strm0_data_valid  ;

  input                                         std__mgr39__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane20_strm1_data        ;
  output                                        mgr39__std__lane20_strm1_data_valid  ;

  input                                         std__mgr39__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane21_strm0_data        ;
  output                                        mgr39__std__lane21_strm0_data_valid  ;

  input                                         std__mgr39__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane21_strm1_data        ;
  output                                        mgr39__std__lane21_strm1_data_valid  ;

  input                                         std__mgr39__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane22_strm0_data        ;
  output                                        mgr39__std__lane22_strm0_data_valid  ;

  input                                         std__mgr39__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane22_strm1_data        ;
  output                                        mgr39__std__lane22_strm1_data_valid  ;

  input                                         std__mgr39__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane23_strm0_data        ;
  output                                        mgr39__std__lane23_strm0_data_valid  ;

  input                                         std__mgr39__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane23_strm1_data        ;
  output                                        mgr39__std__lane23_strm1_data_valid  ;

  input                                         std__mgr39__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane24_strm0_data        ;
  output                                        mgr39__std__lane24_strm0_data_valid  ;

  input                                         std__mgr39__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane24_strm1_data        ;
  output                                        mgr39__std__lane24_strm1_data_valid  ;

  input                                         std__mgr39__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane25_strm0_data        ;
  output                                        mgr39__std__lane25_strm0_data_valid  ;

  input                                         std__mgr39__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane25_strm1_data        ;
  output                                        mgr39__std__lane25_strm1_data_valid  ;

  input                                         std__mgr39__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane26_strm0_data        ;
  output                                        mgr39__std__lane26_strm0_data_valid  ;

  input                                         std__mgr39__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane26_strm1_data        ;
  output                                        mgr39__std__lane26_strm1_data_valid  ;

  input                                         std__mgr39__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane27_strm0_data        ;
  output                                        mgr39__std__lane27_strm0_data_valid  ;

  input                                         std__mgr39__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane27_strm1_data        ;
  output                                        mgr39__std__lane27_strm1_data_valid  ;

  input                                         std__mgr39__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane28_strm0_data        ;
  output                                        mgr39__std__lane28_strm0_data_valid  ;

  input                                         std__mgr39__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane28_strm1_data        ;
  output                                        mgr39__std__lane28_strm1_data_valid  ;

  input                                         std__mgr39__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane29_strm0_data        ;
  output                                        mgr39__std__lane29_strm0_data_valid  ;

  input                                         std__mgr39__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane29_strm1_data        ;
  output                                        mgr39__std__lane29_strm1_data_valid  ;

  input                                         std__mgr39__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane30_strm0_data        ;
  output                                        mgr39__std__lane30_strm0_data_valid  ;

  input                                         std__mgr39__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane30_strm1_data        ;
  output                                        mgr39__std__lane30_strm1_data_valid  ;

  input                                         std__mgr39__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane31_strm0_data        ;
  output                                        mgr39__std__lane31_strm0_data_valid  ;

  input                                         std__mgr39__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane31_strm1_data        ;
  output                                        mgr39__std__lane31_strm1_data_valid  ;

  input                                         std__mgr40__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane0_strm0_data        ;
  output                                        mgr40__std__lane0_strm0_data_valid  ;

  input                                         std__mgr40__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane0_strm1_data        ;
  output                                        mgr40__std__lane0_strm1_data_valid  ;

  input                                         std__mgr40__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane1_strm0_data        ;
  output                                        mgr40__std__lane1_strm0_data_valid  ;

  input                                         std__mgr40__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane1_strm1_data        ;
  output                                        mgr40__std__lane1_strm1_data_valid  ;

  input                                         std__mgr40__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane2_strm0_data        ;
  output                                        mgr40__std__lane2_strm0_data_valid  ;

  input                                         std__mgr40__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane2_strm1_data        ;
  output                                        mgr40__std__lane2_strm1_data_valid  ;

  input                                         std__mgr40__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane3_strm0_data        ;
  output                                        mgr40__std__lane3_strm0_data_valid  ;

  input                                         std__mgr40__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane3_strm1_data        ;
  output                                        mgr40__std__lane3_strm1_data_valid  ;

  input                                         std__mgr40__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane4_strm0_data        ;
  output                                        mgr40__std__lane4_strm0_data_valid  ;

  input                                         std__mgr40__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane4_strm1_data        ;
  output                                        mgr40__std__lane4_strm1_data_valid  ;

  input                                         std__mgr40__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane5_strm0_data        ;
  output                                        mgr40__std__lane5_strm0_data_valid  ;

  input                                         std__mgr40__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane5_strm1_data        ;
  output                                        mgr40__std__lane5_strm1_data_valid  ;

  input                                         std__mgr40__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane6_strm0_data        ;
  output                                        mgr40__std__lane6_strm0_data_valid  ;

  input                                         std__mgr40__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane6_strm1_data        ;
  output                                        mgr40__std__lane6_strm1_data_valid  ;

  input                                         std__mgr40__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane7_strm0_data        ;
  output                                        mgr40__std__lane7_strm0_data_valid  ;

  input                                         std__mgr40__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane7_strm1_data        ;
  output                                        mgr40__std__lane7_strm1_data_valid  ;

  input                                         std__mgr40__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane8_strm0_data        ;
  output                                        mgr40__std__lane8_strm0_data_valid  ;

  input                                         std__mgr40__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane8_strm1_data        ;
  output                                        mgr40__std__lane8_strm1_data_valid  ;

  input                                         std__mgr40__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane9_strm0_data        ;
  output                                        mgr40__std__lane9_strm0_data_valid  ;

  input                                         std__mgr40__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane9_strm1_data        ;
  output                                        mgr40__std__lane9_strm1_data_valid  ;

  input                                         std__mgr40__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane10_strm0_data        ;
  output                                        mgr40__std__lane10_strm0_data_valid  ;

  input                                         std__mgr40__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane10_strm1_data        ;
  output                                        mgr40__std__lane10_strm1_data_valid  ;

  input                                         std__mgr40__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane11_strm0_data        ;
  output                                        mgr40__std__lane11_strm0_data_valid  ;

  input                                         std__mgr40__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane11_strm1_data        ;
  output                                        mgr40__std__lane11_strm1_data_valid  ;

  input                                         std__mgr40__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane12_strm0_data        ;
  output                                        mgr40__std__lane12_strm0_data_valid  ;

  input                                         std__mgr40__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane12_strm1_data        ;
  output                                        mgr40__std__lane12_strm1_data_valid  ;

  input                                         std__mgr40__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane13_strm0_data        ;
  output                                        mgr40__std__lane13_strm0_data_valid  ;

  input                                         std__mgr40__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane13_strm1_data        ;
  output                                        mgr40__std__lane13_strm1_data_valid  ;

  input                                         std__mgr40__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane14_strm0_data        ;
  output                                        mgr40__std__lane14_strm0_data_valid  ;

  input                                         std__mgr40__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane14_strm1_data        ;
  output                                        mgr40__std__lane14_strm1_data_valid  ;

  input                                         std__mgr40__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane15_strm0_data        ;
  output                                        mgr40__std__lane15_strm0_data_valid  ;

  input                                         std__mgr40__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane15_strm1_data        ;
  output                                        mgr40__std__lane15_strm1_data_valid  ;

  input                                         std__mgr40__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane16_strm0_data        ;
  output                                        mgr40__std__lane16_strm0_data_valid  ;

  input                                         std__mgr40__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane16_strm1_data        ;
  output                                        mgr40__std__lane16_strm1_data_valid  ;

  input                                         std__mgr40__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane17_strm0_data        ;
  output                                        mgr40__std__lane17_strm0_data_valid  ;

  input                                         std__mgr40__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane17_strm1_data        ;
  output                                        mgr40__std__lane17_strm1_data_valid  ;

  input                                         std__mgr40__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane18_strm0_data        ;
  output                                        mgr40__std__lane18_strm0_data_valid  ;

  input                                         std__mgr40__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane18_strm1_data        ;
  output                                        mgr40__std__lane18_strm1_data_valid  ;

  input                                         std__mgr40__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane19_strm0_data        ;
  output                                        mgr40__std__lane19_strm0_data_valid  ;

  input                                         std__mgr40__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane19_strm1_data        ;
  output                                        mgr40__std__lane19_strm1_data_valid  ;

  input                                         std__mgr40__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane20_strm0_data        ;
  output                                        mgr40__std__lane20_strm0_data_valid  ;

  input                                         std__mgr40__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane20_strm1_data        ;
  output                                        mgr40__std__lane20_strm1_data_valid  ;

  input                                         std__mgr40__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane21_strm0_data        ;
  output                                        mgr40__std__lane21_strm0_data_valid  ;

  input                                         std__mgr40__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane21_strm1_data        ;
  output                                        mgr40__std__lane21_strm1_data_valid  ;

  input                                         std__mgr40__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane22_strm0_data        ;
  output                                        mgr40__std__lane22_strm0_data_valid  ;

  input                                         std__mgr40__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane22_strm1_data        ;
  output                                        mgr40__std__lane22_strm1_data_valid  ;

  input                                         std__mgr40__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane23_strm0_data        ;
  output                                        mgr40__std__lane23_strm0_data_valid  ;

  input                                         std__mgr40__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane23_strm1_data        ;
  output                                        mgr40__std__lane23_strm1_data_valid  ;

  input                                         std__mgr40__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane24_strm0_data        ;
  output                                        mgr40__std__lane24_strm0_data_valid  ;

  input                                         std__mgr40__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane24_strm1_data        ;
  output                                        mgr40__std__lane24_strm1_data_valid  ;

  input                                         std__mgr40__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane25_strm0_data        ;
  output                                        mgr40__std__lane25_strm0_data_valid  ;

  input                                         std__mgr40__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane25_strm1_data        ;
  output                                        mgr40__std__lane25_strm1_data_valid  ;

  input                                         std__mgr40__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane26_strm0_data        ;
  output                                        mgr40__std__lane26_strm0_data_valid  ;

  input                                         std__mgr40__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane26_strm1_data        ;
  output                                        mgr40__std__lane26_strm1_data_valid  ;

  input                                         std__mgr40__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane27_strm0_data        ;
  output                                        mgr40__std__lane27_strm0_data_valid  ;

  input                                         std__mgr40__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane27_strm1_data        ;
  output                                        mgr40__std__lane27_strm1_data_valid  ;

  input                                         std__mgr40__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane28_strm0_data        ;
  output                                        mgr40__std__lane28_strm0_data_valid  ;

  input                                         std__mgr40__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane28_strm1_data        ;
  output                                        mgr40__std__lane28_strm1_data_valid  ;

  input                                         std__mgr40__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane29_strm0_data        ;
  output                                        mgr40__std__lane29_strm0_data_valid  ;

  input                                         std__mgr40__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane29_strm1_data        ;
  output                                        mgr40__std__lane29_strm1_data_valid  ;

  input                                         std__mgr40__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane30_strm0_data        ;
  output                                        mgr40__std__lane30_strm0_data_valid  ;

  input                                         std__mgr40__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane30_strm1_data        ;
  output                                        mgr40__std__lane30_strm1_data_valid  ;

  input                                         std__mgr40__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane31_strm0_data        ;
  output                                        mgr40__std__lane31_strm0_data_valid  ;

  input                                         std__mgr40__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane31_strm1_data        ;
  output                                        mgr40__std__lane31_strm1_data_valid  ;

  input                                         std__mgr41__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane0_strm0_data        ;
  output                                        mgr41__std__lane0_strm0_data_valid  ;

  input                                         std__mgr41__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane0_strm1_data        ;
  output                                        mgr41__std__lane0_strm1_data_valid  ;

  input                                         std__mgr41__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane1_strm0_data        ;
  output                                        mgr41__std__lane1_strm0_data_valid  ;

  input                                         std__mgr41__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane1_strm1_data        ;
  output                                        mgr41__std__lane1_strm1_data_valid  ;

  input                                         std__mgr41__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane2_strm0_data        ;
  output                                        mgr41__std__lane2_strm0_data_valid  ;

  input                                         std__mgr41__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane2_strm1_data        ;
  output                                        mgr41__std__lane2_strm1_data_valid  ;

  input                                         std__mgr41__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane3_strm0_data        ;
  output                                        mgr41__std__lane3_strm0_data_valid  ;

  input                                         std__mgr41__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane3_strm1_data        ;
  output                                        mgr41__std__lane3_strm1_data_valid  ;

  input                                         std__mgr41__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane4_strm0_data        ;
  output                                        mgr41__std__lane4_strm0_data_valid  ;

  input                                         std__mgr41__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane4_strm1_data        ;
  output                                        mgr41__std__lane4_strm1_data_valid  ;

  input                                         std__mgr41__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane5_strm0_data        ;
  output                                        mgr41__std__lane5_strm0_data_valid  ;

  input                                         std__mgr41__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane5_strm1_data        ;
  output                                        mgr41__std__lane5_strm1_data_valid  ;

  input                                         std__mgr41__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane6_strm0_data        ;
  output                                        mgr41__std__lane6_strm0_data_valid  ;

  input                                         std__mgr41__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane6_strm1_data        ;
  output                                        mgr41__std__lane6_strm1_data_valid  ;

  input                                         std__mgr41__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane7_strm0_data        ;
  output                                        mgr41__std__lane7_strm0_data_valid  ;

  input                                         std__mgr41__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane7_strm1_data        ;
  output                                        mgr41__std__lane7_strm1_data_valid  ;

  input                                         std__mgr41__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane8_strm0_data        ;
  output                                        mgr41__std__lane8_strm0_data_valid  ;

  input                                         std__mgr41__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane8_strm1_data        ;
  output                                        mgr41__std__lane8_strm1_data_valid  ;

  input                                         std__mgr41__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane9_strm0_data        ;
  output                                        mgr41__std__lane9_strm0_data_valid  ;

  input                                         std__mgr41__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane9_strm1_data        ;
  output                                        mgr41__std__lane9_strm1_data_valid  ;

  input                                         std__mgr41__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane10_strm0_data        ;
  output                                        mgr41__std__lane10_strm0_data_valid  ;

  input                                         std__mgr41__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane10_strm1_data        ;
  output                                        mgr41__std__lane10_strm1_data_valid  ;

  input                                         std__mgr41__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane11_strm0_data        ;
  output                                        mgr41__std__lane11_strm0_data_valid  ;

  input                                         std__mgr41__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane11_strm1_data        ;
  output                                        mgr41__std__lane11_strm1_data_valid  ;

  input                                         std__mgr41__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane12_strm0_data        ;
  output                                        mgr41__std__lane12_strm0_data_valid  ;

  input                                         std__mgr41__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane12_strm1_data        ;
  output                                        mgr41__std__lane12_strm1_data_valid  ;

  input                                         std__mgr41__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane13_strm0_data        ;
  output                                        mgr41__std__lane13_strm0_data_valid  ;

  input                                         std__mgr41__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane13_strm1_data        ;
  output                                        mgr41__std__lane13_strm1_data_valid  ;

  input                                         std__mgr41__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane14_strm0_data        ;
  output                                        mgr41__std__lane14_strm0_data_valid  ;

  input                                         std__mgr41__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane14_strm1_data        ;
  output                                        mgr41__std__lane14_strm1_data_valid  ;

  input                                         std__mgr41__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane15_strm0_data        ;
  output                                        mgr41__std__lane15_strm0_data_valid  ;

  input                                         std__mgr41__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane15_strm1_data        ;
  output                                        mgr41__std__lane15_strm1_data_valid  ;

  input                                         std__mgr41__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane16_strm0_data        ;
  output                                        mgr41__std__lane16_strm0_data_valid  ;

  input                                         std__mgr41__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane16_strm1_data        ;
  output                                        mgr41__std__lane16_strm1_data_valid  ;

  input                                         std__mgr41__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane17_strm0_data        ;
  output                                        mgr41__std__lane17_strm0_data_valid  ;

  input                                         std__mgr41__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane17_strm1_data        ;
  output                                        mgr41__std__lane17_strm1_data_valid  ;

  input                                         std__mgr41__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane18_strm0_data        ;
  output                                        mgr41__std__lane18_strm0_data_valid  ;

  input                                         std__mgr41__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane18_strm1_data        ;
  output                                        mgr41__std__lane18_strm1_data_valid  ;

  input                                         std__mgr41__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane19_strm0_data        ;
  output                                        mgr41__std__lane19_strm0_data_valid  ;

  input                                         std__mgr41__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane19_strm1_data        ;
  output                                        mgr41__std__lane19_strm1_data_valid  ;

  input                                         std__mgr41__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane20_strm0_data        ;
  output                                        mgr41__std__lane20_strm0_data_valid  ;

  input                                         std__mgr41__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane20_strm1_data        ;
  output                                        mgr41__std__lane20_strm1_data_valid  ;

  input                                         std__mgr41__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane21_strm0_data        ;
  output                                        mgr41__std__lane21_strm0_data_valid  ;

  input                                         std__mgr41__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane21_strm1_data        ;
  output                                        mgr41__std__lane21_strm1_data_valid  ;

  input                                         std__mgr41__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane22_strm0_data        ;
  output                                        mgr41__std__lane22_strm0_data_valid  ;

  input                                         std__mgr41__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane22_strm1_data        ;
  output                                        mgr41__std__lane22_strm1_data_valid  ;

  input                                         std__mgr41__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane23_strm0_data        ;
  output                                        mgr41__std__lane23_strm0_data_valid  ;

  input                                         std__mgr41__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane23_strm1_data        ;
  output                                        mgr41__std__lane23_strm1_data_valid  ;

  input                                         std__mgr41__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane24_strm0_data        ;
  output                                        mgr41__std__lane24_strm0_data_valid  ;

  input                                         std__mgr41__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane24_strm1_data        ;
  output                                        mgr41__std__lane24_strm1_data_valid  ;

  input                                         std__mgr41__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane25_strm0_data        ;
  output                                        mgr41__std__lane25_strm0_data_valid  ;

  input                                         std__mgr41__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane25_strm1_data        ;
  output                                        mgr41__std__lane25_strm1_data_valid  ;

  input                                         std__mgr41__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane26_strm0_data        ;
  output                                        mgr41__std__lane26_strm0_data_valid  ;

  input                                         std__mgr41__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane26_strm1_data        ;
  output                                        mgr41__std__lane26_strm1_data_valid  ;

  input                                         std__mgr41__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane27_strm0_data        ;
  output                                        mgr41__std__lane27_strm0_data_valid  ;

  input                                         std__mgr41__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane27_strm1_data        ;
  output                                        mgr41__std__lane27_strm1_data_valid  ;

  input                                         std__mgr41__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane28_strm0_data        ;
  output                                        mgr41__std__lane28_strm0_data_valid  ;

  input                                         std__mgr41__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane28_strm1_data        ;
  output                                        mgr41__std__lane28_strm1_data_valid  ;

  input                                         std__mgr41__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane29_strm0_data        ;
  output                                        mgr41__std__lane29_strm0_data_valid  ;

  input                                         std__mgr41__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane29_strm1_data        ;
  output                                        mgr41__std__lane29_strm1_data_valid  ;

  input                                         std__mgr41__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane30_strm0_data        ;
  output                                        mgr41__std__lane30_strm0_data_valid  ;

  input                                         std__mgr41__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane30_strm1_data        ;
  output                                        mgr41__std__lane30_strm1_data_valid  ;

  input                                         std__mgr41__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane31_strm0_data        ;
  output                                        mgr41__std__lane31_strm0_data_valid  ;

  input                                         std__mgr41__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane31_strm1_data        ;
  output                                        mgr41__std__lane31_strm1_data_valid  ;

  input                                         std__mgr42__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane0_strm0_data        ;
  output                                        mgr42__std__lane0_strm0_data_valid  ;

  input                                         std__mgr42__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane0_strm1_data        ;
  output                                        mgr42__std__lane0_strm1_data_valid  ;

  input                                         std__mgr42__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane1_strm0_data        ;
  output                                        mgr42__std__lane1_strm0_data_valid  ;

  input                                         std__mgr42__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane1_strm1_data        ;
  output                                        mgr42__std__lane1_strm1_data_valid  ;

  input                                         std__mgr42__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane2_strm0_data        ;
  output                                        mgr42__std__lane2_strm0_data_valid  ;

  input                                         std__mgr42__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane2_strm1_data        ;
  output                                        mgr42__std__lane2_strm1_data_valid  ;

  input                                         std__mgr42__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane3_strm0_data        ;
  output                                        mgr42__std__lane3_strm0_data_valid  ;

  input                                         std__mgr42__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane3_strm1_data        ;
  output                                        mgr42__std__lane3_strm1_data_valid  ;

  input                                         std__mgr42__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane4_strm0_data        ;
  output                                        mgr42__std__lane4_strm0_data_valid  ;

  input                                         std__mgr42__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane4_strm1_data        ;
  output                                        mgr42__std__lane4_strm1_data_valid  ;

  input                                         std__mgr42__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane5_strm0_data        ;
  output                                        mgr42__std__lane5_strm0_data_valid  ;

  input                                         std__mgr42__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane5_strm1_data        ;
  output                                        mgr42__std__lane5_strm1_data_valid  ;

  input                                         std__mgr42__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane6_strm0_data        ;
  output                                        mgr42__std__lane6_strm0_data_valid  ;

  input                                         std__mgr42__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane6_strm1_data        ;
  output                                        mgr42__std__lane6_strm1_data_valid  ;

  input                                         std__mgr42__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane7_strm0_data        ;
  output                                        mgr42__std__lane7_strm0_data_valid  ;

  input                                         std__mgr42__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane7_strm1_data        ;
  output                                        mgr42__std__lane7_strm1_data_valid  ;

  input                                         std__mgr42__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane8_strm0_data        ;
  output                                        mgr42__std__lane8_strm0_data_valid  ;

  input                                         std__mgr42__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane8_strm1_data        ;
  output                                        mgr42__std__lane8_strm1_data_valid  ;

  input                                         std__mgr42__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane9_strm0_data        ;
  output                                        mgr42__std__lane9_strm0_data_valid  ;

  input                                         std__mgr42__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane9_strm1_data        ;
  output                                        mgr42__std__lane9_strm1_data_valid  ;

  input                                         std__mgr42__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane10_strm0_data        ;
  output                                        mgr42__std__lane10_strm0_data_valid  ;

  input                                         std__mgr42__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane10_strm1_data        ;
  output                                        mgr42__std__lane10_strm1_data_valid  ;

  input                                         std__mgr42__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane11_strm0_data        ;
  output                                        mgr42__std__lane11_strm0_data_valid  ;

  input                                         std__mgr42__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane11_strm1_data        ;
  output                                        mgr42__std__lane11_strm1_data_valid  ;

  input                                         std__mgr42__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane12_strm0_data        ;
  output                                        mgr42__std__lane12_strm0_data_valid  ;

  input                                         std__mgr42__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane12_strm1_data        ;
  output                                        mgr42__std__lane12_strm1_data_valid  ;

  input                                         std__mgr42__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane13_strm0_data        ;
  output                                        mgr42__std__lane13_strm0_data_valid  ;

  input                                         std__mgr42__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane13_strm1_data        ;
  output                                        mgr42__std__lane13_strm1_data_valid  ;

  input                                         std__mgr42__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane14_strm0_data        ;
  output                                        mgr42__std__lane14_strm0_data_valid  ;

  input                                         std__mgr42__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane14_strm1_data        ;
  output                                        mgr42__std__lane14_strm1_data_valid  ;

  input                                         std__mgr42__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane15_strm0_data        ;
  output                                        mgr42__std__lane15_strm0_data_valid  ;

  input                                         std__mgr42__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane15_strm1_data        ;
  output                                        mgr42__std__lane15_strm1_data_valid  ;

  input                                         std__mgr42__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane16_strm0_data        ;
  output                                        mgr42__std__lane16_strm0_data_valid  ;

  input                                         std__mgr42__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane16_strm1_data        ;
  output                                        mgr42__std__lane16_strm1_data_valid  ;

  input                                         std__mgr42__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane17_strm0_data        ;
  output                                        mgr42__std__lane17_strm0_data_valid  ;

  input                                         std__mgr42__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane17_strm1_data        ;
  output                                        mgr42__std__lane17_strm1_data_valid  ;

  input                                         std__mgr42__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane18_strm0_data        ;
  output                                        mgr42__std__lane18_strm0_data_valid  ;

  input                                         std__mgr42__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane18_strm1_data        ;
  output                                        mgr42__std__lane18_strm1_data_valid  ;

  input                                         std__mgr42__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane19_strm0_data        ;
  output                                        mgr42__std__lane19_strm0_data_valid  ;

  input                                         std__mgr42__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane19_strm1_data        ;
  output                                        mgr42__std__lane19_strm1_data_valid  ;

  input                                         std__mgr42__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane20_strm0_data        ;
  output                                        mgr42__std__lane20_strm0_data_valid  ;

  input                                         std__mgr42__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane20_strm1_data        ;
  output                                        mgr42__std__lane20_strm1_data_valid  ;

  input                                         std__mgr42__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane21_strm0_data        ;
  output                                        mgr42__std__lane21_strm0_data_valid  ;

  input                                         std__mgr42__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane21_strm1_data        ;
  output                                        mgr42__std__lane21_strm1_data_valid  ;

  input                                         std__mgr42__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane22_strm0_data        ;
  output                                        mgr42__std__lane22_strm0_data_valid  ;

  input                                         std__mgr42__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane22_strm1_data        ;
  output                                        mgr42__std__lane22_strm1_data_valid  ;

  input                                         std__mgr42__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane23_strm0_data        ;
  output                                        mgr42__std__lane23_strm0_data_valid  ;

  input                                         std__mgr42__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane23_strm1_data        ;
  output                                        mgr42__std__lane23_strm1_data_valid  ;

  input                                         std__mgr42__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane24_strm0_data        ;
  output                                        mgr42__std__lane24_strm0_data_valid  ;

  input                                         std__mgr42__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane24_strm1_data        ;
  output                                        mgr42__std__lane24_strm1_data_valid  ;

  input                                         std__mgr42__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane25_strm0_data        ;
  output                                        mgr42__std__lane25_strm0_data_valid  ;

  input                                         std__mgr42__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane25_strm1_data        ;
  output                                        mgr42__std__lane25_strm1_data_valid  ;

  input                                         std__mgr42__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane26_strm0_data        ;
  output                                        mgr42__std__lane26_strm0_data_valid  ;

  input                                         std__mgr42__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane26_strm1_data        ;
  output                                        mgr42__std__lane26_strm1_data_valid  ;

  input                                         std__mgr42__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane27_strm0_data        ;
  output                                        mgr42__std__lane27_strm0_data_valid  ;

  input                                         std__mgr42__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane27_strm1_data        ;
  output                                        mgr42__std__lane27_strm1_data_valid  ;

  input                                         std__mgr42__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane28_strm0_data        ;
  output                                        mgr42__std__lane28_strm0_data_valid  ;

  input                                         std__mgr42__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane28_strm1_data        ;
  output                                        mgr42__std__lane28_strm1_data_valid  ;

  input                                         std__mgr42__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane29_strm0_data        ;
  output                                        mgr42__std__lane29_strm0_data_valid  ;

  input                                         std__mgr42__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane29_strm1_data        ;
  output                                        mgr42__std__lane29_strm1_data_valid  ;

  input                                         std__mgr42__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane30_strm0_data        ;
  output                                        mgr42__std__lane30_strm0_data_valid  ;

  input                                         std__mgr42__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane30_strm1_data        ;
  output                                        mgr42__std__lane30_strm1_data_valid  ;

  input                                         std__mgr42__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane31_strm0_data        ;
  output                                        mgr42__std__lane31_strm0_data_valid  ;

  input                                         std__mgr42__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane31_strm1_data        ;
  output                                        mgr42__std__lane31_strm1_data_valid  ;

  input                                         std__mgr43__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane0_strm0_data        ;
  output                                        mgr43__std__lane0_strm0_data_valid  ;

  input                                         std__mgr43__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane0_strm1_data        ;
  output                                        mgr43__std__lane0_strm1_data_valid  ;

  input                                         std__mgr43__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane1_strm0_data        ;
  output                                        mgr43__std__lane1_strm0_data_valid  ;

  input                                         std__mgr43__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane1_strm1_data        ;
  output                                        mgr43__std__lane1_strm1_data_valid  ;

  input                                         std__mgr43__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane2_strm0_data        ;
  output                                        mgr43__std__lane2_strm0_data_valid  ;

  input                                         std__mgr43__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane2_strm1_data        ;
  output                                        mgr43__std__lane2_strm1_data_valid  ;

  input                                         std__mgr43__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane3_strm0_data        ;
  output                                        mgr43__std__lane3_strm0_data_valid  ;

  input                                         std__mgr43__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane3_strm1_data        ;
  output                                        mgr43__std__lane3_strm1_data_valid  ;

  input                                         std__mgr43__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane4_strm0_data        ;
  output                                        mgr43__std__lane4_strm0_data_valid  ;

  input                                         std__mgr43__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane4_strm1_data        ;
  output                                        mgr43__std__lane4_strm1_data_valid  ;

  input                                         std__mgr43__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane5_strm0_data        ;
  output                                        mgr43__std__lane5_strm0_data_valid  ;

  input                                         std__mgr43__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane5_strm1_data        ;
  output                                        mgr43__std__lane5_strm1_data_valid  ;

  input                                         std__mgr43__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane6_strm0_data        ;
  output                                        mgr43__std__lane6_strm0_data_valid  ;

  input                                         std__mgr43__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane6_strm1_data        ;
  output                                        mgr43__std__lane6_strm1_data_valid  ;

  input                                         std__mgr43__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane7_strm0_data        ;
  output                                        mgr43__std__lane7_strm0_data_valid  ;

  input                                         std__mgr43__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane7_strm1_data        ;
  output                                        mgr43__std__lane7_strm1_data_valid  ;

  input                                         std__mgr43__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane8_strm0_data        ;
  output                                        mgr43__std__lane8_strm0_data_valid  ;

  input                                         std__mgr43__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane8_strm1_data        ;
  output                                        mgr43__std__lane8_strm1_data_valid  ;

  input                                         std__mgr43__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane9_strm0_data        ;
  output                                        mgr43__std__lane9_strm0_data_valid  ;

  input                                         std__mgr43__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane9_strm1_data        ;
  output                                        mgr43__std__lane9_strm1_data_valid  ;

  input                                         std__mgr43__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane10_strm0_data        ;
  output                                        mgr43__std__lane10_strm0_data_valid  ;

  input                                         std__mgr43__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane10_strm1_data        ;
  output                                        mgr43__std__lane10_strm1_data_valid  ;

  input                                         std__mgr43__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane11_strm0_data        ;
  output                                        mgr43__std__lane11_strm0_data_valid  ;

  input                                         std__mgr43__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane11_strm1_data        ;
  output                                        mgr43__std__lane11_strm1_data_valid  ;

  input                                         std__mgr43__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane12_strm0_data        ;
  output                                        mgr43__std__lane12_strm0_data_valid  ;

  input                                         std__mgr43__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane12_strm1_data        ;
  output                                        mgr43__std__lane12_strm1_data_valid  ;

  input                                         std__mgr43__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane13_strm0_data        ;
  output                                        mgr43__std__lane13_strm0_data_valid  ;

  input                                         std__mgr43__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane13_strm1_data        ;
  output                                        mgr43__std__lane13_strm1_data_valid  ;

  input                                         std__mgr43__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane14_strm0_data        ;
  output                                        mgr43__std__lane14_strm0_data_valid  ;

  input                                         std__mgr43__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane14_strm1_data        ;
  output                                        mgr43__std__lane14_strm1_data_valid  ;

  input                                         std__mgr43__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane15_strm0_data        ;
  output                                        mgr43__std__lane15_strm0_data_valid  ;

  input                                         std__mgr43__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane15_strm1_data        ;
  output                                        mgr43__std__lane15_strm1_data_valid  ;

  input                                         std__mgr43__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane16_strm0_data        ;
  output                                        mgr43__std__lane16_strm0_data_valid  ;

  input                                         std__mgr43__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane16_strm1_data        ;
  output                                        mgr43__std__lane16_strm1_data_valid  ;

  input                                         std__mgr43__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane17_strm0_data        ;
  output                                        mgr43__std__lane17_strm0_data_valid  ;

  input                                         std__mgr43__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane17_strm1_data        ;
  output                                        mgr43__std__lane17_strm1_data_valid  ;

  input                                         std__mgr43__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane18_strm0_data        ;
  output                                        mgr43__std__lane18_strm0_data_valid  ;

  input                                         std__mgr43__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane18_strm1_data        ;
  output                                        mgr43__std__lane18_strm1_data_valid  ;

  input                                         std__mgr43__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane19_strm0_data        ;
  output                                        mgr43__std__lane19_strm0_data_valid  ;

  input                                         std__mgr43__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane19_strm1_data        ;
  output                                        mgr43__std__lane19_strm1_data_valid  ;

  input                                         std__mgr43__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane20_strm0_data        ;
  output                                        mgr43__std__lane20_strm0_data_valid  ;

  input                                         std__mgr43__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane20_strm1_data        ;
  output                                        mgr43__std__lane20_strm1_data_valid  ;

  input                                         std__mgr43__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane21_strm0_data        ;
  output                                        mgr43__std__lane21_strm0_data_valid  ;

  input                                         std__mgr43__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane21_strm1_data        ;
  output                                        mgr43__std__lane21_strm1_data_valid  ;

  input                                         std__mgr43__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane22_strm0_data        ;
  output                                        mgr43__std__lane22_strm0_data_valid  ;

  input                                         std__mgr43__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane22_strm1_data        ;
  output                                        mgr43__std__lane22_strm1_data_valid  ;

  input                                         std__mgr43__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane23_strm0_data        ;
  output                                        mgr43__std__lane23_strm0_data_valid  ;

  input                                         std__mgr43__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane23_strm1_data        ;
  output                                        mgr43__std__lane23_strm1_data_valid  ;

  input                                         std__mgr43__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane24_strm0_data        ;
  output                                        mgr43__std__lane24_strm0_data_valid  ;

  input                                         std__mgr43__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane24_strm1_data        ;
  output                                        mgr43__std__lane24_strm1_data_valid  ;

  input                                         std__mgr43__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane25_strm0_data        ;
  output                                        mgr43__std__lane25_strm0_data_valid  ;

  input                                         std__mgr43__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane25_strm1_data        ;
  output                                        mgr43__std__lane25_strm1_data_valid  ;

  input                                         std__mgr43__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane26_strm0_data        ;
  output                                        mgr43__std__lane26_strm0_data_valid  ;

  input                                         std__mgr43__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane26_strm1_data        ;
  output                                        mgr43__std__lane26_strm1_data_valid  ;

  input                                         std__mgr43__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane27_strm0_data        ;
  output                                        mgr43__std__lane27_strm0_data_valid  ;

  input                                         std__mgr43__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane27_strm1_data        ;
  output                                        mgr43__std__lane27_strm1_data_valid  ;

  input                                         std__mgr43__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane28_strm0_data        ;
  output                                        mgr43__std__lane28_strm0_data_valid  ;

  input                                         std__mgr43__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane28_strm1_data        ;
  output                                        mgr43__std__lane28_strm1_data_valid  ;

  input                                         std__mgr43__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane29_strm0_data        ;
  output                                        mgr43__std__lane29_strm0_data_valid  ;

  input                                         std__mgr43__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane29_strm1_data        ;
  output                                        mgr43__std__lane29_strm1_data_valid  ;

  input                                         std__mgr43__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane30_strm0_data        ;
  output                                        mgr43__std__lane30_strm0_data_valid  ;

  input                                         std__mgr43__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane30_strm1_data        ;
  output                                        mgr43__std__lane30_strm1_data_valid  ;

  input                                         std__mgr43__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane31_strm0_data        ;
  output                                        mgr43__std__lane31_strm0_data_valid  ;

  input                                         std__mgr43__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane31_strm1_data        ;
  output                                        mgr43__std__lane31_strm1_data_valid  ;

  input                                         std__mgr44__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane0_strm0_data        ;
  output                                        mgr44__std__lane0_strm0_data_valid  ;

  input                                         std__mgr44__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane0_strm1_data        ;
  output                                        mgr44__std__lane0_strm1_data_valid  ;

  input                                         std__mgr44__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane1_strm0_data        ;
  output                                        mgr44__std__lane1_strm0_data_valid  ;

  input                                         std__mgr44__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane1_strm1_data        ;
  output                                        mgr44__std__lane1_strm1_data_valid  ;

  input                                         std__mgr44__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane2_strm0_data        ;
  output                                        mgr44__std__lane2_strm0_data_valid  ;

  input                                         std__mgr44__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane2_strm1_data        ;
  output                                        mgr44__std__lane2_strm1_data_valid  ;

  input                                         std__mgr44__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane3_strm0_data        ;
  output                                        mgr44__std__lane3_strm0_data_valid  ;

  input                                         std__mgr44__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane3_strm1_data        ;
  output                                        mgr44__std__lane3_strm1_data_valid  ;

  input                                         std__mgr44__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane4_strm0_data        ;
  output                                        mgr44__std__lane4_strm0_data_valid  ;

  input                                         std__mgr44__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane4_strm1_data        ;
  output                                        mgr44__std__lane4_strm1_data_valid  ;

  input                                         std__mgr44__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane5_strm0_data        ;
  output                                        mgr44__std__lane5_strm0_data_valid  ;

  input                                         std__mgr44__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane5_strm1_data        ;
  output                                        mgr44__std__lane5_strm1_data_valid  ;

  input                                         std__mgr44__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane6_strm0_data        ;
  output                                        mgr44__std__lane6_strm0_data_valid  ;

  input                                         std__mgr44__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane6_strm1_data        ;
  output                                        mgr44__std__lane6_strm1_data_valid  ;

  input                                         std__mgr44__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane7_strm0_data        ;
  output                                        mgr44__std__lane7_strm0_data_valid  ;

  input                                         std__mgr44__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane7_strm1_data        ;
  output                                        mgr44__std__lane7_strm1_data_valid  ;

  input                                         std__mgr44__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane8_strm0_data        ;
  output                                        mgr44__std__lane8_strm0_data_valid  ;

  input                                         std__mgr44__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane8_strm1_data        ;
  output                                        mgr44__std__lane8_strm1_data_valid  ;

  input                                         std__mgr44__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane9_strm0_data        ;
  output                                        mgr44__std__lane9_strm0_data_valid  ;

  input                                         std__mgr44__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane9_strm1_data        ;
  output                                        mgr44__std__lane9_strm1_data_valid  ;

  input                                         std__mgr44__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane10_strm0_data        ;
  output                                        mgr44__std__lane10_strm0_data_valid  ;

  input                                         std__mgr44__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane10_strm1_data        ;
  output                                        mgr44__std__lane10_strm1_data_valid  ;

  input                                         std__mgr44__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane11_strm0_data        ;
  output                                        mgr44__std__lane11_strm0_data_valid  ;

  input                                         std__mgr44__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane11_strm1_data        ;
  output                                        mgr44__std__lane11_strm1_data_valid  ;

  input                                         std__mgr44__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane12_strm0_data        ;
  output                                        mgr44__std__lane12_strm0_data_valid  ;

  input                                         std__mgr44__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane12_strm1_data        ;
  output                                        mgr44__std__lane12_strm1_data_valid  ;

  input                                         std__mgr44__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane13_strm0_data        ;
  output                                        mgr44__std__lane13_strm0_data_valid  ;

  input                                         std__mgr44__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane13_strm1_data        ;
  output                                        mgr44__std__lane13_strm1_data_valid  ;

  input                                         std__mgr44__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane14_strm0_data        ;
  output                                        mgr44__std__lane14_strm0_data_valid  ;

  input                                         std__mgr44__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane14_strm1_data        ;
  output                                        mgr44__std__lane14_strm1_data_valid  ;

  input                                         std__mgr44__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane15_strm0_data        ;
  output                                        mgr44__std__lane15_strm0_data_valid  ;

  input                                         std__mgr44__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane15_strm1_data        ;
  output                                        mgr44__std__lane15_strm1_data_valid  ;

  input                                         std__mgr44__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane16_strm0_data        ;
  output                                        mgr44__std__lane16_strm0_data_valid  ;

  input                                         std__mgr44__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane16_strm1_data        ;
  output                                        mgr44__std__lane16_strm1_data_valid  ;

  input                                         std__mgr44__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane17_strm0_data        ;
  output                                        mgr44__std__lane17_strm0_data_valid  ;

  input                                         std__mgr44__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane17_strm1_data        ;
  output                                        mgr44__std__lane17_strm1_data_valid  ;

  input                                         std__mgr44__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane18_strm0_data        ;
  output                                        mgr44__std__lane18_strm0_data_valid  ;

  input                                         std__mgr44__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane18_strm1_data        ;
  output                                        mgr44__std__lane18_strm1_data_valid  ;

  input                                         std__mgr44__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane19_strm0_data        ;
  output                                        mgr44__std__lane19_strm0_data_valid  ;

  input                                         std__mgr44__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane19_strm1_data        ;
  output                                        mgr44__std__lane19_strm1_data_valid  ;

  input                                         std__mgr44__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane20_strm0_data        ;
  output                                        mgr44__std__lane20_strm0_data_valid  ;

  input                                         std__mgr44__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane20_strm1_data        ;
  output                                        mgr44__std__lane20_strm1_data_valid  ;

  input                                         std__mgr44__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane21_strm0_data        ;
  output                                        mgr44__std__lane21_strm0_data_valid  ;

  input                                         std__mgr44__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane21_strm1_data        ;
  output                                        mgr44__std__lane21_strm1_data_valid  ;

  input                                         std__mgr44__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane22_strm0_data        ;
  output                                        mgr44__std__lane22_strm0_data_valid  ;

  input                                         std__mgr44__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane22_strm1_data        ;
  output                                        mgr44__std__lane22_strm1_data_valid  ;

  input                                         std__mgr44__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane23_strm0_data        ;
  output                                        mgr44__std__lane23_strm0_data_valid  ;

  input                                         std__mgr44__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane23_strm1_data        ;
  output                                        mgr44__std__lane23_strm1_data_valid  ;

  input                                         std__mgr44__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane24_strm0_data        ;
  output                                        mgr44__std__lane24_strm0_data_valid  ;

  input                                         std__mgr44__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane24_strm1_data        ;
  output                                        mgr44__std__lane24_strm1_data_valid  ;

  input                                         std__mgr44__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane25_strm0_data        ;
  output                                        mgr44__std__lane25_strm0_data_valid  ;

  input                                         std__mgr44__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane25_strm1_data        ;
  output                                        mgr44__std__lane25_strm1_data_valid  ;

  input                                         std__mgr44__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane26_strm0_data        ;
  output                                        mgr44__std__lane26_strm0_data_valid  ;

  input                                         std__mgr44__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane26_strm1_data        ;
  output                                        mgr44__std__lane26_strm1_data_valid  ;

  input                                         std__mgr44__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane27_strm0_data        ;
  output                                        mgr44__std__lane27_strm0_data_valid  ;

  input                                         std__mgr44__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane27_strm1_data        ;
  output                                        mgr44__std__lane27_strm1_data_valid  ;

  input                                         std__mgr44__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane28_strm0_data        ;
  output                                        mgr44__std__lane28_strm0_data_valid  ;

  input                                         std__mgr44__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane28_strm1_data        ;
  output                                        mgr44__std__lane28_strm1_data_valid  ;

  input                                         std__mgr44__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane29_strm0_data        ;
  output                                        mgr44__std__lane29_strm0_data_valid  ;

  input                                         std__mgr44__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane29_strm1_data        ;
  output                                        mgr44__std__lane29_strm1_data_valid  ;

  input                                         std__mgr44__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane30_strm0_data        ;
  output                                        mgr44__std__lane30_strm0_data_valid  ;

  input                                         std__mgr44__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane30_strm1_data        ;
  output                                        mgr44__std__lane30_strm1_data_valid  ;

  input                                         std__mgr44__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane31_strm0_data        ;
  output                                        mgr44__std__lane31_strm0_data_valid  ;

  input                                         std__mgr44__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane31_strm1_data        ;
  output                                        mgr44__std__lane31_strm1_data_valid  ;

  input                                         std__mgr45__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane0_strm0_data        ;
  output                                        mgr45__std__lane0_strm0_data_valid  ;

  input                                         std__mgr45__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane0_strm1_data        ;
  output                                        mgr45__std__lane0_strm1_data_valid  ;

  input                                         std__mgr45__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane1_strm0_data        ;
  output                                        mgr45__std__lane1_strm0_data_valid  ;

  input                                         std__mgr45__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane1_strm1_data        ;
  output                                        mgr45__std__lane1_strm1_data_valid  ;

  input                                         std__mgr45__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane2_strm0_data        ;
  output                                        mgr45__std__lane2_strm0_data_valid  ;

  input                                         std__mgr45__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane2_strm1_data        ;
  output                                        mgr45__std__lane2_strm1_data_valid  ;

  input                                         std__mgr45__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane3_strm0_data        ;
  output                                        mgr45__std__lane3_strm0_data_valid  ;

  input                                         std__mgr45__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane3_strm1_data        ;
  output                                        mgr45__std__lane3_strm1_data_valid  ;

  input                                         std__mgr45__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane4_strm0_data        ;
  output                                        mgr45__std__lane4_strm0_data_valid  ;

  input                                         std__mgr45__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane4_strm1_data        ;
  output                                        mgr45__std__lane4_strm1_data_valid  ;

  input                                         std__mgr45__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane5_strm0_data        ;
  output                                        mgr45__std__lane5_strm0_data_valid  ;

  input                                         std__mgr45__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane5_strm1_data        ;
  output                                        mgr45__std__lane5_strm1_data_valid  ;

  input                                         std__mgr45__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane6_strm0_data        ;
  output                                        mgr45__std__lane6_strm0_data_valid  ;

  input                                         std__mgr45__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane6_strm1_data        ;
  output                                        mgr45__std__lane6_strm1_data_valid  ;

  input                                         std__mgr45__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane7_strm0_data        ;
  output                                        mgr45__std__lane7_strm0_data_valid  ;

  input                                         std__mgr45__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane7_strm1_data        ;
  output                                        mgr45__std__lane7_strm1_data_valid  ;

  input                                         std__mgr45__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane8_strm0_data        ;
  output                                        mgr45__std__lane8_strm0_data_valid  ;

  input                                         std__mgr45__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane8_strm1_data        ;
  output                                        mgr45__std__lane8_strm1_data_valid  ;

  input                                         std__mgr45__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane9_strm0_data        ;
  output                                        mgr45__std__lane9_strm0_data_valid  ;

  input                                         std__mgr45__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane9_strm1_data        ;
  output                                        mgr45__std__lane9_strm1_data_valid  ;

  input                                         std__mgr45__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane10_strm0_data        ;
  output                                        mgr45__std__lane10_strm0_data_valid  ;

  input                                         std__mgr45__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane10_strm1_data        ;
  output                                        mgr45__std__lane10_strm1_data_valid  ;

  input                                         std__mgr45__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane11_strm0_data        ;
  output                                        mgr45__std__lane11_strm0_data_valid  ;

  input                                         std__mgr45__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane11_strm1_data        ;
  output                                        mgr45__std__lane11_strm1_data_valid  ;

  input                                         std__mgr45__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane12_strm0_data        ;
  output                                        mgr45__std__lane12_strm0_data_valid  ;

  input                                         std__mgr45__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane12_strm1_data        ;
  output                                        mgr45__std__lane12_strm1_data_valid  ;

  input                                         std__mgr45__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane13_strm0_data        ;
  output                                        mgr45__std__lane13_strm0_data_valid  ;

  input                                         std__mgr45__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane13_strm1_data        ;
  output                                        mgr45__std__lane13_strm1_data_valid  ;

  input                                         std__mgr45__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane14_strm0_data        ;
  output                                        mgr45__std__lane14_strm0_data_valid  ;

  input                                         std__mgr45__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane14_strm1_data        ;
  output                                        mgr45__std__lane14_strm1_data_valid  ;

  input                                         std__mgr45__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane15_strm0_data        ;
  output                                        mgr45__std__lane15_strm0_data_valid  ;

  input                                         std__mgr45__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane15_strm1_data        ;
  output                                        mgr45__std__lane15_strm1_data_valid  ;

  input                                         std__mgr45__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane16_strm0_data        ;
  output                                        mgr45__std__lane16_strm0_data_valid  ;

  input                                         std__mgr45__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane16_strm1_data        ;
  output                                        mgr45__std__lane16_strm1_data_valid  ;

  input                                         std__mgr45__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane17_strm0_data        ;
  output                                        mgr45__std__lane17_strm0_data_valid  ;

  input                                         std__mgr45__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane17_strm1_data        ;
  output                                        mgr45__std__lane17_strm1_data_valid  ;

  input                                         std__mgr45__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane18_strm0_data        ;
  output                                        mgr45__std__lane18_strm0_data_valid  ;

  input                                         std__mgr45__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane18_strm1_data        ;
  output                                        mgr45__std__lane18_strm1_data_valid  ;

  input                                         std__mgr45__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane19_strm0_data        ;
  output                                        mgr45__std__lane19_strm0_data_valid  ;

  input                                         std__mgr45__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane19_strm1_data        ;
  output                                        mgr45__std__lane19_strm1_data_valid  ;

  input                                         std__mgr45__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane20_strm0_data        ;
  output                                        mgr45__std__lane20_strm0_data_valid  ;

  input                                         std__mgr45__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane20_strm1_data        ;
  output                                        mgr45__std__lane20_strm1_data_valid  ;

  input                                         std__mgr45__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane21_strm0_data        ;
  output                                        mgr45__std__lane21_strm0_data_valid  ;

  input                                         std__mgr45__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane21_strm1_data        ;
  output                                        mgr45__std__lane21_strm1_data_valid  ;

  input                                         std__mgr45__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane22_strm0_data        ;
  output                                        mgr45__std__lane22_strm0_data_valid  ;

  input                                         std__mgr45__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane22_strm1_data        ;
  output                                        mgr45__std__lane22_strm1_data_valid  ;

  input                                         std__mgr45__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane23_strm0_data        ;
  output                                        mgr45__std__lane23_strm0_data_valid  ;

  input                                         std__mgr45__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane23_strm1_data        ;
  output                                        mgr45__std__lane23_strm1_data_valid  ;

  input                                         std__mgr45__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane24_strm0_data        ;
  output                                        mgr45__std__lane24_strm0_data_valid  ;

  input                                         std__mgr45__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane24_strm1_data        ;
  output                                        mgr45__std__lane24_strm1_data_valid  ;

  input                                         std__mgr45__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane25_strm0_data        ;
  output                                        mgr45__std__lane25_strm0_data_valid  ;

  input                                         std__mgr45__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane25_strm1_data        ;
  output                                        mgr45__std__lane25_strm1_data_valid  ;

  input                                         std__mgr45__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane26_strm0_data        ;
  output                                        mgr45__std__lane26_strm0_data_valid  ;

  input                                         std__mgr45__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane26_strm1_data        ;
  output                                        mgr45__std__lane26_strm1_data_valid  ;

  input                                         std__mgr45__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane27_strm0_data        ;
  output                                        mgr45__std__lane27_strm0_data_valid  ;

  input                                         std__mgr45__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane27_strm1_data        ;
  output                                        mgr45__std__lane27_strm1_data_valid  ;

  input                                         std__mgr45__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane28_strm0_data        ;
  output                                        mgr45__std__lane28_strm0_data_valid  ;

  input                                         std__mgr45__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane28_strm1_data        ;
  output                                        mgr45__std__lane28_strm1_data_valid  ;

  input                                         std__mgr45__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane29_strm0_data        ;
  output                                        mgr45__std__lane29_strm0_data_valid  ;

  input                                         std__mgr45__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane29_strm1_data        ;
  output                                        mgr45__std__lane29_strm1_data_valid  ;

  input                                         std__mgr45__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane30_strm0_data        ;
  output                                        mgr45__std__lane30_strm0_data_valid  ;

  input                                         std__mgr45__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane30_strm1_data        ;
  output                                        mgr45__std__lane30_strm1_data_valid  ;

  input                                         std__mgr45__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane31_strm0_data        ;
  output                                        mgr45__std__lane31_strm0_data_valid  ;

  input                                         std__mgr45__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane31_strm1_data        ;
  output                                        mgr45__std__lane31_strm1_data_valid  ;

  input                                         std__mgr46__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane0_strm0_data        ;
  output                                        mgr46__std__lane0_strm0_data_valid  ;

  input                                         std__mgr46__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane0_strm1_data        ;
  output                                        mgr46__std__lane0_strm1_data_valid  ;

  input                                         std__mgr46__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane1_strm0_data        ;
  output                                        mgr46__std__lane1_strm0_data_valid  ;

  input                                         std__mgr46__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane1_strm1_data        ;
  output                                        mgr46__std__lane1_strm1_data_valid  ;

  input                                         std__mgr46__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane2_strm0_data        ;
  output                                        mgr46__std__lane2_strm0_data_valid  ;

  input                                         std__mgr46__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane2_strm1_data        ;
  output                                        mgr46__std__lane2_strm1_data_valid  ;

  input                                         std__mgr46__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane3_strm0_data        ;
  output                                        mgr46__std__lane3_strm0_data_valid  ;

  input                                         std__mgr46__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane3_strm1_data        ;
  output                                        mgr46__std__lane3_strm1_data_valid  ;

  input                                         std__mgr46__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane4_strm0_data        ;
  output                                        mgr46__std__lane4_strm0_data_valid  ;

  input                                         std__mgr46__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane4_strm1_data        ;
  output                                        mgr46__std__lane4_strm1_data_valid  ;

  input                                         std__mgr46__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane5_strm0_data        ;
  output                                        mgr46__std__lane5_strm0_data_valid  ;

  input                                         std__mgr46__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane5_strm1_data        ;
  output                                        mgr46__std__lane5_strm1_data_valid  ;

  input                                         std__mgr46__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane6_strm0_data        ;
  output                                        mgr46__std__lane6_strm0_data_valid  ;

  input                                         std__mgr46__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane6_strm1_data        ;
  output                                        mgr46__std__lane6_strm1_data_valid  ;

  input                                         std__mgr46__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane7_strm0_data        ;
  output                                        mgr46__std__lane7_strm0_data_valid  ;

  input                                         std__mgr46__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane7_strm1_data        ;
  output                                        mgr46__std__lane7_strm1_data_valid  ;

  input                                         std__mgr46__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane8_strm0_data        ;
  output                                        mgr46__std__lane8_strm0_data_valid  ;

  input                                         std__mgr46__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane8_strm1_data        ;
  output                                        mgr46__std__lane8_strm1_data_valid  ;

  input                                         std__mgr46__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane9_strm0_data        ;
  output                                        mgr46__std__lane9_strm0_data_valid  ;

  input                                         std__mgr46__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane9_strm1_data        ;
  output                                        mgr46__std__lane9_strm1_data_valid  ;

  input                                         std__mgr46__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane10_strm0_data        ;
  output                                        mgr46__std__lane10_strm0_data_valid  ;

  input                                         std__mgr46__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane10_strm1_data        ;
  output                                        mgr46__std__lane10_strm1_data_valid  ;

  input                                         std__mgr46__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane11_strm0_data        ;
  output                                        mgr46__std__lane11_strm0_data_valid  ;

  input                                         std__mgr46__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane11_strm1_data        ;
  output                                        mgr46__std__lane11_strm1_data_valid  ;

  input                                         std__mgr46__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane12_strm0_data        ;
  output                                        mgr46__std__lane12_strm0_data_valid  ;

  input                                         std__mgr46__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane12_strm1_data        ;
  output                                        mgr46__std__lane12_strm1_data_valid  ;

  input                                         std__mgr46__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane13_strm0_data        ;
  output                                        mgr46__std__lane13_strm0_data_valid  ;

  input                                         std__mgr46__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane13_strm1_data        ;
  output                                        mgr46__std__lane13_strm1_data_valid  ;

  input                                         std__mgr46__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane14_strm0_data        ;
  output                                        mgr46__std__lane14_strm0_data_valid  ;

  input                                         std__mgr46__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane14_strm1_data        ;
  output                                        mgr46__std__lane14_strm1_data_valid  ;

  input                                         std__mgr46__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane15_strm0_data        ;
  output                                        mgr46__std__lane15_strm0_data_valid  ;

  input                                         std__mgr46__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane15_strm1_data        ;
  output                                        mgr46__std__lane15_strm1_data_valid  ;

  input                                         std__mgr46__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane16_strm0_data        ;
  output                                        mgr46__std__lane16_strm0_data_valid  ;

  input                                         std__mgr46__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane16_strm1_data        ;
  output                                        mgr46__std__lane16_strm1_data_valid  ;

  input                                         std__mgr46__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane17_strm0_data        ;
  output                                        mgr46__std__lane17_strm0_data_valid  ;

  input                                         std__mgr46__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane17_strm1_data        ;
  output                                        mgr46__std__lane17_strm1_data_valid  ;

  input                                         std__mgr46__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane18_strm0_data        ;
  output                                        mgr46__std__lane18_strm0_data_valid  ;

  input                                         std__mgr46__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane18_strm1_data        ;
  output                                        mgr46__std__lane18_strm1_data_valid  ;

  input                                         std__mgr46__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane19_strm0_data        ;
  output                                        mgr46__std__lane19_strm0_data_valid  ;

  input                                         std__mgr46__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane19_strm1_data        ;
  output                                        mgr46__std__lane19_strm1_data_valid  ;

  input                                         std__mgr46__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane20_strm0_data        ;
  output                                        mgr46__std__lane20_strm0_data_valid  ;

  input                                         std__mgr46__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane20_strm1_data        ;
  output                                        mgr46__std__lane20_strm1_data_valid  ;

  input                                         std__mgr46__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane21_strm0_data        ;
  output                                        mgr46__std__lane21_strm0_data_valid  ;

  input                                         std__mgr46__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane21_strm1_data        ;
  output                                        mgr46__std__lane21_strm1_data_valid  ;

  input                                         std__mgr46__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane22_strm0_data        ;
  output                                        mgr46__std__lane22_strm0_data_valid  ;

  input                                         std__mgr46__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane22_strm1_data        ;
  output                                        mgr46__std__lane22_strm1_data_valid  ;

  input                                         std__mgr46__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane23_strm0_data        ;
  output                                        mgr46__std__lane23_strm0_data_valid  ;

  input                                         std__mgr46__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane23_strm1_data        ;
  output                                        mgr46__std__lane23_strm1_data_valid  ;

  input                                         std__mgr46__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane24_strm0_data        ;
  output                                        mgr46__std__lane24_strm0_data_valid  ;

  input                                         std__mgr46__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane24_strm1_data        ;
  output                                        mgr46__std__lane24_strm1_data_valid  ;

  input                                         std__mgr46__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane25_strm0_data        ;
  output                                        mgr46__std__lane25_strm0_data_valid  ;

  input                                         std__mgr46__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane25_strm1_data        ;
  output                                        mgr46__std__lane25_strm1_data_valid  ;

  input                                         std__mgr46__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane26_strm0_data        ;
  output                                        mgr46__std__lane26_strm0_data_valid  ;

  input                                         std__mgr46__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane26_strm1_data        ;
  output                                        mgr46__std__lane26_strm1_data_valid  ;

  input                                         std__mgr46__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane27_strm0_data        ;
  output                                        mgr46__std__lane27_strm0_data_valid  ;

  input                                         std__mgr46__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane27_strm1_data        ;
  output                                        mgr46__std__lane27_strm1_data_valid  ;

  input                                         std__mgr46__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane28_strm0_data        ;
  output                                        mgr46__std__lane28_strm0_data_valid  ;

  input                                         std__mgr46__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane28_strm1_data        ;
  output                                        mgr46__std__lane28_strm1_data_valid  ;

  input                                         std__mgr46__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane29_strm0_data        ;
  output                                        mgr46__std__lane29_strm0_data_valid  ;

  input                                         std__mgr46__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane29_strm1_data        ;
  output                                        mgr46__std__lane29_strm1_data_valid  ;

  input                                         std__mgr46__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane30_strm0_data        ;
  output                                        mgr46__std__lane30_strm0_data_valid  ;

  input                                         std__mgr46__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane30_strm1_data        ;
  output                                        mgr46__std__lane30_strm1_data_valid  ;

  input                                         std__mgr46__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane31_strm0_data        ;
  output                                        mgr46__std__lane31_strm0_data_valid  ;

  input                                         std__mgr46__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane31_strm1_data        ;
  output                                        mgr46__std__lane31_strm1_data_valid  ;

  input                                         std__mgr47__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane0_strm0_data        ;
  output                                        mgr47__std__lane0_strm0_data_valid  ;

  input                                         std__mgr47__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane0_strm1_data        ;
  output                                        mgr47__std__lane0_strm1_data_valid  ;

  input                                         std__mgr47__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane1_strm0_data        ;
  output                                        mgr47__std__lane1_strm0_data_valid  ;

  input                                         std__mgr47__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane1_strm1_data        ;
  output                                        mgr47__std__lane1_strm1_data_valid  ;

  input                                         std__mgr47__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane2_strm0_data        ;
  output                                        mgr47__std__lane2_strm0_data_valid  ;

  input                                         std__mgr47__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane2_strm1_data        ;
  output                                        mgr47__std__lane2_strm1_data_valid  ;

  input                                         std__mgr47__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane3_strm0_data        ;
  output                                        mgr47__std__lane3_strm0_data_valid  ;

  input                                         std__mgr47__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane3_strm1_data        ;
  output                                        mgr47__std__lane3_strm1_data_valid  ;

  input                                         std__mgr47__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane4_strm0_data        ;
  output                                        mgr47__std__lane4_strm0_data_valid  ;

  input                                         std__mgr47__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane4_strm1_data        ;
  output                                        mgr47__std__lane4_strm1_data_valid  ;

  input                                         std__mgr47__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane5_strm0_data        ;
  output                                        mgr47__std__lane5_strm0_data_valid  ;

  input                                         std__mgr47__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane5_strm1_data        ;
  output                                        mgr47__std__lane5_strm1_data_valid  ;

  input                                         std__mgr47__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane6_strm0_data        ;
  output                                        mgr47__std__lane6_strm0_data_valid  ;

  input                                         std__mgr47__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane6_strm1_data        ;
  output                                        mgr47__std__lane6_strm1_data_valid  ;

  input                                         std__mgr47__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane7_strm0_data        ;
  output                                        mgr47__std__lane7_strm0_data_valid  ;

  input                                         std__mgr47__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane7_strm1_data        ;
  output                                        mgr47__std__lane7_strm1_data_valid  ;

  input                                         std__mgr47__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane8_strm0_data        ;
  output                                        mgr47__std__lane8_strm0_data_valid  ;

  input                                         std__mgr47__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane8_strm1_data        ;
  output                                        mgr47__std__lane8_strm1_data_valid  ;

  input                                         std__mgr47__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane9_strm0_data        ;
  output                                        mgr47__std__lane9_strm0_data_valid  ;

  input                                         std__mgr47__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane9_strm1_data        ;
  output                                        mgr47__std__lane9_strm1_data_valid  ;

  input                                         std__mgr47__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane10_strm0_data        ;
  output                                        mgr47__std__lane10_strm0_data_valid  ;

  input                                         std__mgr47__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane10_strm1_data        ;
  output                                        mgr47__std__lane10_strm1_data_valid  ;

  input                                         std__mgr47__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane11_strm0_data        ;
  output                                        mgr47__std__lane11_strm0_data_valid  ;

  input                                         std__mgr47__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane11_strm1_data        ;
  output                                        mgr47__std__lane11_strm1_data_valid  ;

  input                                         std__mgr47__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane12_strm0_data        ;
  output                                        mgr47__std__lane12_strm0_data_valid  ;

  input                                         std__mgr47__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane12_strm1_data        ;
  output                                        mgr47__std__lane12_strm1_data_valid  ;

  input                                         std__mgr47__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane13_strm0_data        ;
  output                                        mgr47__std__lane13_strm0_data_valid  ;

  input                                         std__mgr47__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane13_strm1_data        ;
  output                                        mgr47__std__lane13_strm1_data_valid  ;

  input                                         std__mgr47__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane14_strm0_data        ;
  output                                        mgr47__std__lane14_strm0_data_valid  ;

  input                                         std__mgr47__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane14_strm1_data        ;
  output                                        mgr47__std__lane14_strm1_data_valid  ;

  input                                         std__mgr47__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane15_strm0_data        ;
  output                                        mgr47__std__lane15_strm0_data_valid  ;

  input                                         std__mgr47__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane15_strm1_data        ;
  output                                        mgr47__std__lane15_strm1_data_valid  ;

  input                                         std__mgr47__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane16_strm0_data        ;
  output                                        mgr47__std__lane16_strm0_data_valid  ;

  input                                         std__mgr47__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane16_strm1_data        ;
  output                                        mgr47__std__lane16_strm1_data_valid  ;

  input                                         std__mgr47__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane17_strm0_data        ;
  output                                        mgr47__std__lane17_strm0_data_valid  ;

  input                                         std__mgr47__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane17_strm1_data        ;
  output                                        mgr47__std__lane17_strm1_data_valid  ;

  input                                         std__mgr47__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane18_strm0_data        ;
  output                                        mgr47__std__lane18_strm0_data_valid  ;

  input                                         std__mgr47__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane18_strm1_data        ;
  output                                        mgr47__std__lane18_strm1_data_valid  ;

  input                                         std__mgr47__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane19_strm0_data        ;
  output                                        mgr47__std__lane19_strm0_data_valid  ;

  input                                         std__mgr47__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane19_strm1_data        ;
  output                                        mgr47__std__lane19_strm1_data_valid  ;

  input                                         std__mgr47__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane20_strm0_data        ;
  output                                        mgr47__std__lane20_strm0_data_valid  ;

  input                                         std__mgr47__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane20_strm1_data        ;
  output                                        mgr47__std__lane20_strm1_data_valid  ;

  input                                         std__mgr47__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane21_strm0_data        ;
  output                                        mgr47__std__lane21_strm0_data_valid  ;

  input                                         std__mgr47__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane21_strm1_data        ;
  output                                        mgr47__std__lane21_strm1_data_valid  ;

  input                                         std__mgr47__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane22_strm0_data        ;
  output                                        mgr47__std__lane22_strm0_data_valid  ;

  input                                         std__mgr47__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane22_strm1_data        ;
  output                                        mgr47__std__lane22_strm1_data_valid  ;

  input                                         std__mgr47__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane23_strm0_data        ;
  output                                        mgr47__std__lane23_strm0_data_valid  ;

  input                                         std__mgr47__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane23_strm1_data        ;
  output                                        mgr47__std__lane23_strm1_data_valid  ;

  input                                         std__mgr47__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane24_strm0_data        ;
  output                                        mgr47__std__lane24_strm0_data_valid  ;

  input                                         std__mgr47__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane24_strm1_data        ;
  output                                        mgr47__std__lane24_strm1_data_valid  ;

  input                                         std__mgr47__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane25_strm0_data        ;
  output                                        mgr47__std__lane25_strm0_data_valid  ;

  input                                         std__mgr47__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane25_strm1_data        ;
  output                                        mgr47__std__lane25_strm1_data_valid  ;

  input                                         std__mgr47__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane26_strm0_data        ;
  output                                        mgr47__std__lane26_strm0_data_valid  ;

  input                                         std__mgr47__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane26_strm1_data        ;
  output                                        mgr47__std__lane26_strm1_data_valid  ;

  input                                         std__mgr47__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane27_strm0_data        ;
  output                                        mgr47__std__lane27_strm0_data_valid  ;

  input                                         std__mgr47__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane27_strm1_data        ;
  output                                        mgr47__std__lane27_strm1_data_valid  ;

  input                                         std__mgr47__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane28_strm0_data        ;
  output                                        mgr47__std__lane28_strm0_data_valid  ;

  input                                         std__mgr47__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane28_strm1_data        ;
  output                                        mgr47__std__lane28_strm1_data_valid  ;

  input                                         std__mgr47__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane29_strm0_data        ;
  output                                        mgr47__std__lane29_strm0_data_valid  ;

  input                                         std__mgr47__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane29_strm1_data        ;
  output                                        mgr47__std__lane29_strm1_data_valid  ;

  input                                         std__mgr47__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane30_strm0_data        ;
  output                                        mgr47__std__lane30_strm0_data_valid  ;

  input                                         std__mgr47__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane30_strm1_data        ;
  output                                        mgr47__std__lane30_strm1_data_valid  ;

  input                                         std__mgr47__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane31_strm0_data        ;
  output                                        mgr47__std__lane31_strm0_data_valid  ;

  input                                         std__mgr47__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane31_strm1_data        ;
  output                                        mgr47__std__lane31_strm1_data_valid  ;

  input                                         std__mgr48__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane0_strm0_data        ;
  output                                        mgr48__std__lane0_strm0_data_valid  ;

  input                                         std__mgr48__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane0_strm1_data        ;
  output                                        mgr48__std__lane0_strm1_data_valid  ;

  input                                         std__mgr48__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane1_strm0_data        ;
  output                                        mgr48__std__lane1_strm0_data_valid  ;

  input                                         std__mgr48__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane1_strm1_data        ;
  output                                        mgr48__std__lane1_strm1_data_valid  ;

  input                                         std__mgr48__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane2_strm0_data        ;
  output                                        mgr48__std__lane2_strm0_data_valid  ;

  input                                         std__mgr48__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane2_strm1_data        ;
  output                                        mgr48__std__lane2_strm1_data_valid  ;

  input                                         std__mgr48__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane3_strm0_data        ;
  output                                        mgr48__std__lane3_strm0_data_valid  ;

  input                                         std__mgr48__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane3_strm1_data        ;
  output                                        mgr48__std__lane3_strm1_data_valid  ;

  input                                         std__mgr48__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane4_strm0_data        ;
  output                                        mgr48__std__lane4_strm0_data_valid  ;

  input                                         std__mgr48__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane4_strm1_data        ;
  output                                        mgr48__std__lane4_strm1_data_valid  ;

  input                                         std__mgr48__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane5_strm0_data        ;
  output                                        mgr48__std__lane5_strm0_data_valid  ;

  input                                         std__mgr48__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane5_strm1_data        ;
  output                                        mgr48__std__lane5_strm1_data_valid  ;

  input                                         std__mgr48__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane6_strm0_data        ;
  output                                        mgr48__std__lane6_strm0_data_valid  ;

  input                                         std__mgr48__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane6_strm1_data        ;
  output                                        mgr48__std__lane6_strm1_data_valid  ;

  input                                         std__mgr48__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane7_strm0_data        ;
  output                                        mgr48__std__lane7_strm0_data_valid  ;

  input                                         std__mgr48__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane7_strm1_data        ;
  output                                        mgr48__std__lane7_strm1_data_valid  ;

  input                                         std__mgr48__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane8_strm0_data        ;
  output                                        mgr48__std__lane8_strm0_data_valid  ;

  input                                         std__mgr48__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane8_strm1_data        ;
  output                                        mgr48__std__lane8_strm1_data_valid  ;

  input                                         std__mgr48__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane9_strm0_data        ;
  output                                        mgr48__std__lane9_strm0_data_valid  ;

  input                                         std__mgr48__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane9_strm1_data        ;
  output                                        mgr48__std__lane9_strm1_data_valid  ;

  input                                         std__mgr48__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane10_strm0_data        ;
  output                                        mgr48__std__lane10_strm0_data_valid  ;

  input                                         std__mgr48__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane10_strm1_data        ;
  output                                        mgr48__std__lane10_strm1_data_valid  ;

  input                                         std__mgr48__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane11_strm0_data        ;
  output                                        mgr48__std__lane11_strm0_data_valid  ;

  input                                         std__mgr48__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane11_strm1_data        ;
  output                                        mgr48__std__lane11_strm1_data_valid  ;

  input                                         std__mgr48__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane12_strm0_data        ;
  output                                        mgr48__std__lane12_strm0_data_valid  ;

  input                                         std__mgr48__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane12_strm1_data        ;
  output                                        mgr48__std__lane12_strm1_data_valid  ;

  input                                         std__mgr48__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane13_strm0_data        ;
  output                                        mgr48__std__lane13_strm0_data_valid  ;

  input                                         std__mgr48__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane13_strm1_data        ;
  output                                        mgr48__std__lane13_strm1_data_valid  ;

  input                                         std__mgr48__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane14_strm0_data        ;
  output                                        mgr48__std__lane14_strm0_data_valid  ;

  input                                         std__mgr48__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane14_strm1_data        ;
  output                                        mgr48__std__lane14_strm1_data_valid  ;

  input                                         std__mgr48__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane15_strm0_data        ;
  output                                        mgr48__std__lane15_strm0_data_valid  ;

  input                                         std__mgr48__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane15_strm1_data        ;
  output                                        mgr48__std__lane15_strm1_data_valid  ;

  input                                         std__mgr48__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane16_strm0_data        ;
  output                                        mgr48__std__lane16_strm0_data_valid  ;

  input                                         std__mgr48__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane16_strm1_data        ;
  output                                        mgr48__std__lane16_strm1_data_valid  ;

  input                                         std__mgr48__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane17_strm0_data        ;
  output                                        mgr48__std__lane17_strm0_data_valid  ;

  input                                         std__mgr48__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane17_strm1_data        ;
  output                                        mgr48__std__lane17_strm1_data_valid  ;

  input                                         std__mgr48__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane18_strm0_data        ;
  output                                        mgr48__std__lane18_strm0_data_valid  ;

  input                                         std__mgr48__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane18_strm1_data        ;
  output                                        mgr48__std__lane18_strm1_data_valid  ;

  input                                         std__mgr48__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane19_strm0_data        ;
  output                                        mgr48__std__lane19_strm0_data_valid  ;

  input                                         std__mgr48__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane19_strm1_data        ;
  output                                        mgr48__std__lane19_strm1_data_valid  ;

  input                                         std__mgr48__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane20_strm0_data        ;
  output                                        mgr48__std__lane20_strm0_data_valid  ;

  input                                         std__mgr48__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane20_strm1_data        ;
  output                                        mgr48__std__lane20_strm1_data_valid  ;

  input                                         std__mgr48__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane21_strm0_data        ;
  output                                        mgr48__std__lane21_strm0_data_valid  ;

  input                                         std__mgr48__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane21_strm1_data        ;
  output                                        mgr48__std__lane21_strm1_data_valid  ;

  input                                         std__mgr48__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane22_strm0_data        ;
  output                                        mgr48__std__lane22_strm0_data_valid  ;

  input                                         std__mgr48__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane22_strm1_data        ;
  output                                        mgr48__std__lane22_strm1_data_valid  ;

  input                                         std__mgr48__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane23_strm0_data        ;
  output                                        mgr48__std__lane23_strm0_data_valid  ;

  input                                         std__mgr48__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane23_strm1_data        ;
  output                                        mgr48__std__lane23_strm1_data_valid  ;

  input                                         std__mgr48__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane24_strm0_data        ;
  output                                        mgr48__std__lane24_strm0_data_valid  ;

  input                                         std__mgr48__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane24_strm1_data        ;
  output                                        mgr48__std__lane24_strm1_data_valid  ;

  input                                         std__mgr48__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane25_strm0_data        ;
  output                                        mgr48__std__lane25_strm0_data_valid  ;

  input                                         std__mgr48__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane25_strm1_data        ;
  output                                        mgr48__std__lane25_strm1_data_valid  ;

  input                                         std__mgr48__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane26_strm0_data        ;
  output                                        mgr48__std__lane26_strm0_data_valid  ;

  input                                         std__mgr48__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane26_strm1_data        ;
  output                                        mgr48__std__lane26_strm1_data_valid  ;

  input                                         std__mgr48__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane27_strm0_data        ;
  output                                        mgr48__std__lane27_strm0_data_valid  ;

  input                                         std__mgr48__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane27_strm1_data        ;
  output                                        mgr48__std__lane27_strm1_data_valid  ;

  input                                         std__mgr48__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane28_strm0_data        ;
  output                                        mgr48__std__lane28_strm0_data_valid  ;

  input                                         std__mgr48__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane28_strm1_data        ;
  output                                        mgr48__std__lane28_strm1_data_valid  ;

  input                                         std__mgr48__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane29_strm0_data        ;
  output                                        mgr48__std__lane29_strm0_data_valid  ;

  input                                         std__mgr48__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane29_strm1_data        ;
  output                                        mgr48__std__lane29_strm1_data_valid  ;

  input                                         std__mgr48__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane30_strm0_data        ;
  output                                        mgr48__std__lane30_strm0_data_valid  ;

  input                                         std__mgr48__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane30_strm1_data        ;
  output                                        mgr48__std__lane30_strm1_data_valid  ;

  input                                         std__mgr48__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane31_strm0_data        ;
  output                                        mgr48__std__lane31_strm0_data_valid  ;

  input                                         std__mgr48__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane31_strm1_data        ;
  output                                        mgr48__std__lane31_strm1_data_valid  ;

  input                                         std__mgr49__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane0_strm0_data        ;
  output                                        mgr49__std__lane0_strm0_data_valid  ;

  input                                         std__mgr49__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane0_strm1_data        ;
  output                                        mgr49__std__lane0_strm1_data_valid  ;

  input                                         std__mgr49__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane1_strm0_data        ;
  output                                        mgr49__std__lane1_strm0_data_valid  ;

  input                                         std__mgr49__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane1_strm1_data        ;
  output                                        mgr49__std__lane1_strm1_data_valid  ;

  input                                         std__mgr49__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane2_strm0_data        ;
  output                                        mgr49__std__lane2_strm0_data_valid  ;

  input                                         std__mgr49__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane2_strm1_data        ;
  output                                        mgr49__std__lane2_strm1_data_valid  ;

  input                                         std__mgr49__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane3_strm0_data        ;
  output                                        mgr49__std__lane3_strm0_data_valid  ;

  input                                         std__mgr49__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane3_strm1_data        ;
  output                                        mgr49__std__lane3_strm1_data_valid  ;

  input                                         std__mgr49__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane4_strm0_data        ;
  output                                        mgr49__std__lane4_strm0_data_valid  ;

  input                                         std__mgr49__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane4_strm1_data        ;
  output                                        mgr49__std__lane4_strm1_data_valid  ;

  input                                         std__mgr49__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane5_strm0_data        ;
  output                                        mgr49__std__lane5_strm0_data_valid  ;

  input                                         std__mgr49__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane5_strm1_data        ;
  output                                        mgr49__std__lane5_strm1_data_valid  ;

  input                                         std__mgr49__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane6_strm0_data        ;
  output                                        mgr49__std__lane6_strm0_data_valid  ;

  input                                         std__mgr49__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane6_strm1_data        ;
  output                                        mgr49__std__lane6_strm1_data_valid  ;

  input                                         std__mgr49__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane7_strm0_data        ;
  output                                        mgr49__std__lane7_strm0_data_valid  ;

  input                                         std__mgr49__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane7_strm1_data        ;
  output                                        mgr49__std__lane7_strm1_data_valid  ;

  input                                         std__mgr49__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane8_strm0_data        ;
  output                                        mgr49__std__lane8_strm0_data_valid  ;

  input                                         std__mgr49__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane8_strm1_data        ;
  output                                        mgr49__std__lane8_strm1_data_valid  ;

  input                                         std__mgr49__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane9_strm0_data        ;
  output                                        mgr49__std__lane9_strm0_data_valid  ;

  input                                         std__mgr49__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane9_strm1_data        ;
  output                                        mgr49__std__lane9_strm1_data_valid  ;

  input                                         std__mgr49__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane10_strm0_data        ;
  output                                        mgr49__std__lane10_strm0_data_valid  ;

  input                                         std__mgr49__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane10_strm1_data        ;
  output                                        mgr49__std__lane10_strm1_data_valid  ;

  input                                         std__mgr49__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane11_strm0_data        ;
  output                                        mgr49__std__lane11_strm0_data_valid  ;

  input                                         std__mgr49__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane11_strm1_data        ;
  output                                        mgr49__std__lane11_strm1_data_valid  ;

  input                                         std__mgr49__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane12_strm0_data        ;
  output                                        mgr49__std__lane12_strm0_data_valid  ;

  input                                         std__mgr49__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane12_strm1_data        ;
  output                                        mgr49__std__lane12_strm1_data_valid  ;

  input                                         std__mgr49__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane13_strm0_data        ;
  output                                        mgr49__std__lane13_strm0_data_valid  ;

  input                                         std__mgr49__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane13_strm1_data        ;
  output                                        mgr49__std__lane13_strm1_data_valid  ;

  input                                         std__mgr49__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane14_strm0_data        ;
  output                                        mgr49__std__lane14_strm0_data_valid  ;

  input                                         std__mgr49__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane14_strm1_data        ;
  output                                        mgr49__std__lane14_strm1_data_valid  ;

  input                                         std__mgr49__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane15_strm0_data        ;
  output                                        mgr49__std__lane15_strm0_data_valid  ;

  input                                         std__mgr49__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane15_strm1_data        ;
  output                                        mgr49__std__lane15_strm1_data_valid  ;

  input                                         std__mgr49__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane16_strm0_data        ;
  output                                        mgr49__std__lane16_strm0_data_valid  ;

  input                                         std__mgr49__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane16_strm1_data        ;
  output                                        mgr49__std__lane16_strm1_data_valid  ;

  input                                         std__mgr49__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane17_strm0_data        ;
  output                                        mgr49__std__lane17_strm0_data_valid  ;

  input                                         std__mgr49__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane17_strm1_data        ;
  output                                        mgr49__std__lane17_strm1_data_valid  ;

  input                                         std__mgr49__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane18_strm0_data        ;
  output                                        mgr49__std__lane18_strm0_data_valid  ;

  input                                         std__mgr49__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane18_strm1_data        ;
  output                                        mgr49__std__lane18_strm1_data_valid  ;

  input                                         std__mgr49__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane19_strm0_data        ;
  output                                        mgr49__std__lane19_strm0_data_valid  ;

  input                                         std__mgr49__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane19_strm1_data        ;
  output                                        mgr49__std__lane19_strm1_data_valid  ;

  input                                         std__mgr49__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane20_strm0_data        ;
  output                                        mgr49__std__lane20_strm0_data_valid  ;

  input                                         std__mgr49__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane20_strm1_data        ;
  output                                        mgr49__std__lane20_strm1_data_valid  ;

  input                                         std__mgr49__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane21_strm0_data        ;
  output                                        mgr49__std__lane21_strm0_data_valid  ;

  input                                         std__mgr49__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane21_strm1_data        ;
  output                                        mgr49__std__lane21_strm1_data_valid  ;

  input                                         std__mgr49__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane22_strm0_data        ;
  output                                        mgr49__std__lane22_strm0_data_valid  ;

  input                                         std__mgr49__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane22_strm1_data        ;
  output                                        mgr49__std__lane22_strm1_data_valid  ;

  input                                         std__mgr49__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane23_strm0_data        ;
  output                                        mgr49__std__lane23_strm0_data_valid  ;

  input                                         std__mgr49__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane23_strm1_data        ;
  output                                        mgr49__std__lane23_strm1_data_valid  ;

  input                                         std__mgr49__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane24_strm0_data        ;
  output                                        mgr49__std__lane24_strm0_data_valid  ;

  input                                         std__mgr49__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane24_strm1_data        ;
  output                                        mgr49__std__lane24_strm1_data_valid  ;

  input                                         std__mgr49__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane25_strm0_data        ;
  output                                        mgr49__std__lane25_strm0_data_valid  ;

  input                                         std__mgr49__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane25_strm1_data        ;
  output                                        mgr49__std__lane25_strm1_data_valid  ;

  input                                         std__mgr49__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane26_strm0_data        ;
  output                                        mgr49__std__lane26_strm0_data_valid  ;

  input                                         std__mgr49__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane26_strm1_data        ;
  output                                        mgr49__std__lane26_strm1_data_valid  ;

  input                                         std__mgr49__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane27_strm0_data        ;
  output                                        mgr49__std__lane27_strm0_data_valid  ;

  input                                         std__mgr49__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane27_strm1_data        ;
  output                                        mgr49__std__lane27_strm1_data_valid  ;

  input                                         std__mgr49__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane28_strm0_data        ;
  output                                        mgr49__std__lane28_strm0_data_valid  ;

  input                                         std__mgr49__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane28_strm1_data        ;
  output                                        mgr49__std__lane28_strm1_data_valid  ;

  input                                         std__mgr49__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane29_strm0_data        ;
  output                                        mgr49__std__lane29_strm0_data_valid  ;

  input                                         std__mgr49__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane29_strm1_data        ;
  output                                        mgr49__std__lane29_strm1_data_valid  ;

  input                                         std__mgr49__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane30_strm0_data        ;
  output                                        mgr49__std__lane30_strm0_data_valid  ;

  input                                         std__mgr49__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane30_strm1_data        ;
  output                                        mgr49__std__lane30_strm1_data_valid  ;

  input                                         std__mgr49__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane31_strm0_data        ;
  output                                        mgr49__std__lane31_strm0_data_valid  ;

  input                                         std__mgr49__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane31_strm1_data        ;
  output                                        mgr49__std__lane31_strm1_data_valid  ;

  input                                         std__mgr50__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane0_strm0_data        ;
  output                                        mgr50__std__lane0_strm0_data_valid  ;

  input                                         std__mgr50__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane0_strm1_data        ;
  output                                        mgr50__std__lane0_strm1_data_valid  ;

  input                                         std__mgr50__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane1_strm0_data        ;
  output                                        mgr50__std__lane1_strm0_data_valid  ;

  input                                         std__mgr50__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane1_strm1_data        ;
  output                                        mgr50__std__lane1_strm1_data_valid  ;

  input                                         std__mgr50__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane2_strm0_data        ;
  output                                        mgr50__std__lane2_strm0_data_valid  ;

  input                                         std__mgr50__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane2_strm1_data        ;
  output                                        mgr50__std__lane2_strm1_data_valid  ;

  input                                         std__mgr50__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane3_strm0_data        ;
  output                                        mgr50__std__lane3_strm0_data_valid  ;

  input                                         std__mgr50__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane3_strm1_data        ;
  output                                        mgr50__std__lane3_strm1_data_valid  ;

  input                                         std__mgr50__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane4_strm0_data        ;
  output                                        mgr50__std__lane4_strm0_data_valid  ;

  input                                         std__mgr50__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane4_strm1_data        ;
  output                                        mgr50__std__lane4_strm1_data_valid  ;

  input                                         std__mgr50__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane5_strm0_data        ;
  output                                        mgr50__std__lane5_strm0_data_valid  ;

  input                                         std__mgr50__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane5_strm1_data        ;
  output                                        mgr50__std__lane5_strm1_data_valid  ;

  input                                         std__mgr50__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane6_strm0_data        ;
  output                                        mgr50__std__lane6_strm0_data_valid  ;

  input                                         std__mgr50__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane6_strm1_data        ;
  output                                        mgr50__std__lane6_strm1_data_valid  ;

  input                                         std__mgr50__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane7_strm0_data        ;
  output                                        mgr50__std__lane7_strm0_data_valid  ;

  input                                         std__mgr50__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane7_strm1_data        ;
  output                                        mgr50__std__lane7_strm1_data_valid  ;

  input                                         std__mgr50__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane8_strm0_data        ;
  output                                        mgr50__std__lane8_strm0_data_valid  ;

  input                                         std__mgr50__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane8_strm1_data        ;
  output                                        mgr50__std__lane8_strm1_data_valid  ;

  input                                         std__mgr50__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane9_strm0_data        ;
  output                                        mgr50__std__lane9_strm0_data_valid  ;

  input                                         std__mgr50__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane9_strm1_data        ;
  output                                        mgr50__std__lane9_strm1_data_valid  ;

  input                                         std__mgr50__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane10_strm0_data        ;
  output                                        mgr50__std__lane10_strm0_data_valid  ;

  input                                         std__mgr50__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane10_strm1_data        ;
  output                                        mgr50__std__lane10_strm1_data_valid  ;

  input                                         std__mgr50__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane11_strm0_data        ;
  output                                        mgr50__std__lane11_strm0_data_valid  ;

  input                                         std__mgr50__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane11_strm1_data        ;
  output                                        mgr50__std__lane11_strm1_data_valid  ;

  input                                         std__mgr50__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane12_strm0_data        ;
  output                                        mgr50__std__lane12_strm0_data_valid  ;

  input                                         std__mgr50__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane12_strm1_data        ;
  output                                        mgr50__std__lane12_strm1_data_valid  ;

  input                                         std__mgr50__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane13_strm0_data        ;
  output                                        mgr50__std__lane13_strm0_data_valid  ;

  input                                         std__mgr50__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane13_strm1_data        ;
  output                                        mgr50__std__lane13_strm1_data_valid  ;

  input                                         std__mgr50__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane14_strm0_data        ;
  output                                        mgr50__std__lane14_strm0_data_valid  ;

  input                                         std__mgr50__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane14_strm1_data        ;
  output                                        mgr50__std__lane14_strm1_data_valid  ;

  input                                         std__mgr50__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane15_strm0_data        ;
  output                                        mgr50__std__lane15_strm0_data_valid  ;

  input                                         std__mgr50__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane15_strm1_data        ;
  output                                        mgr50__std__lane15_strm1_data_valid  ;

  input                                         std__mgr50__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane16_strm0_data        ;
  output                                        mgr50__std__lane16_strm0_data_valid  ;

  input                                         std__mgr50__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane16_strm1_data        ;
  output                                        mgr50__std__lane16_strm1_data_valid  ;

  input                                         std__mgr50__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane17_strm0_data        ;
  output                                        mgr50__std__lane17_strm0_data_valid  ;

  input                                         std__mgr50__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane17_strm1_data        ;
  output                                        mgr50__std__lane17_strm1_data_valid  ;

  input                                         std__mgr50__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane18_strm0_data        ;
  output                                        mgr50__std__lane18_strm0_data_valid  ;

  input                                         std__mgr50__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane18_strm1_data        ;
  output                                        mgr50__std__lane18_strm1_data_valid  ;

  input                                         std__mgr50__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane19_strm0_data        ;
  output                                        mgr50__std__lane19_strm0_data_valid  ;

  input                                         std__mgr50__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane19_strm1_data        ;
  output                                        mgr50__std__lane19_strm1_data_valid  ;

  input                                         std__mgr50__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane20_strm0_data        ;
  output                                        mgr50__std__lane20_strm0_data_valid  ;

  input                                         std__mgr50__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane20_strm1_data        ;
  output                                        mgr50__std__lane20_strm1_data_valid  ;

  input                                         std__mgr50__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane21_strm0_data        ;
  output                                        mgr50__std__lane21_strm0_data_valid  ;

  input                                         std__mgr50__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane21_strm1_data        ;
  output                                        mgr50__std__lane21_strm1_data_valid  ;

  input                                         std__mgr50__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane22_strm0_data        ;
  output                                        mgr50__std__lane22_strm0_data_valid  ;

  input                                         std__mgr50__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane22_strm1_data        ;
  output                                        mgr50__std__lane22_strm1_data_valid  ;

  input                                         std__mgr50__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane23_strm0_data        ;
  output                                        mgr50__std__lane23_strm0_data_valid  ;

  input                                         std__mgr50__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane23_strm1_data        ;
  output                                        mgr50__std__lane23_strm1_data_valid  ;

  input                                         std__mgr50__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane24_strm0_data        ;
  output                                        mgr50__std__lane24_strm0_data_valid  ;

  input                                         std__mgr50__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane24_strm1_data        ;
  output                                        mgr50__std__lane24_strm1_data_valid  ;

  input                                         std__mgr50__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane25_strm0_data        ;
  output                                        mgr50__std__lane25_strm0_data_valid  ;

  input                                         std__mgr50__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane25_strm1_data        ;
  output                                        mgr50__std__lane25_strm1_data_valid  ;

  input                                         std__mgr50__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane26_strm0_data        ;
  output                                        mgr50__std__lane26_strm0_data_valid  ;

  input                                         std__mgr50__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane26_strm1_data        ;
  output                                        mgr50__std__lane26_strm1_data_valid  ;

  input                                         std__mgr50__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane27_strm0_data        ;
  output                                        mgr50__std__lane27_strm0_data_valid  ;

  input                                         std__mgr50__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane27_strm1_data        ;
  output                                        mgr50__std__lane27_strm1_data_valid  ;

  input                                         std__mgr50__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane28_strm0_data        ;
  output                                        mgr50__std__lane28_strm0_data_valid  ;

  input                                         std__mgr50__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane28_strm1_data        ;
  output                                        mgr50__std__lane28_strm1_data_valid  ;

  input                                         std__mgr50__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane29_strm0_data        ;
  output                                        mgr50__std__lane29_strm0_data_valid  ;

  input                                         std__mgr50__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane29_strm1_data        ;
  output                                        mgr50__std__lane29_strm1_data_valid  ;

  input                                         std__mgr50__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane30_strm0_data        ;
  output                                        mgr50__std__lane30_strm0_data_valid  ;

  input                                         std__mgr50__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane30_strm1_data        ;
  output                                        mgr50__std__lane30_strm1_data_valid  ;

  input                                         std__mgr50__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane31_strm0_data        ;
  output                                        mgr50__std__lane31_strm0_data_valid  ;

  input                                         std__mgr50__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane31_strm1_data        ;
  output                                        mgr50__std__lane31_strm1_data_valid  ;

  input                                         std__mgr51__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane0_strm0_data        ;
  output                                        mgr51__std__lane0_strm0_data_valid  ;

  input                                         std__mgr51__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane0_strm1_data        ;
  output                                        mgr51__std__lane0_strm1_data_valid  ;

  input                                         std__mgr51__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane1_strm0_data        ;
  output                                        mgr51__std__lane1_strm0_data_valid  ;

  input                                         std__mgr51__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane1_strm1_data        ;
  output                                        mgr51__std__lane1_strm1_data_valid  ;

  input                                         std__mgr51__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane2_strm0_data        ;
  output                                        mgr51__std__lane2_strm0_data_valid  ;

  input                                         std__mgr51__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane2_strm1_data        ;
  output                                        mgr51__std__lane2_strm1_data_valid  ;

  input                                         std__mgr51__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane3_strm0_data        ;
  output                                        mgr51__std__lane3_strm0_data_valid  ;

  input                                         std__mgr51__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane3_strm1_data        ;
  output                                        mgr51__std__lane3_strm1_data_valid  ;

  input                                         std__mgr51__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane4_strm0_data        ;
  output                                        mgr51__std__lane4_strm0_data_valid  ;

  input                                         std__mgr51__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane4_strm1_data        ;
  output                                        mgr51__std__lane4_strm1_data_valid  ;

  input                                         std__mgr51__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane5_strm0_data        ;
  output                                        mgr51__std__lane5_strm0_data_valid  ;

  input                                         std__mgr51__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane5_strm1_data        ;
  output                                        mgr51__std__lane5_strm1_data_valid  ;

  input                                         std__mgr51__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane6_strm0_data        ;
  output                                        mgr51__std__lane6_strm0_data_valid  ;

  input                                         std__mgr51__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane6_strm1_data        ;
  output                                        mgr51__std__lane6_strm1_data_valid  ;

  input                                         std__mgr51__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane7_strm0_data        ;
  output                                        mgr51__std__lane7_strm0_data_valid  ;

  input                                         std__mgr51__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane7_strm1_data        ;
  output                                        mgr51__std__lane7_strm1_data_valid  ;

  input                                         std__mgr51__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane8_strm0_data        ;
  output                                        mgr51__std__lane8_strm0_data_valid  ;

  input                                         std__mgr51__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane8_strm1_data        ;
  output                                        mgr51__std__lane8_strm1_data_valid  ;

  input                                         std__mgr51__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane9_strm0_data        ;
  output                                        mgr51__std__lane9_strm0_data_valid  ;

  input                                         std__mgr51__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane9_strm1_data        ;
  output                                        mgr51__std__lane9_strm1_data_valid  ;

  input                                         std__mgr51__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane10_strm0_data        ;
  output                                        mgr51__std__lane10_strm0_data_valid  ;

  input                                         std__mgr51__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane10_strm1_data        ;
  output                                        mgr51__std__lane10_strm1_data_valid  ;

  input                                         std__mgr51__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane11_strm0_data        ;
  output                                        mgr51__std__lane11_strm0_data_valid  ;

  input                                         std__mgr51__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane11_strm1_data        ;
  output                                        mgr51__std__lane11_strm1_data_valid  ;

  input                                         std__mgr51__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane12_strm0_data        ;
  output                                        mgr51__std__lane12_strm0_data_valid  ;

  input                                         std__mgr51__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane12_strm1_data        ;
  output                                        mgr51__std__lane12_strm1_data_valid  ;

  input                                         std__mgr51__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane13_strm0_data        ;
  output                                        mgr51__std__lane13_strm0_data_valid  ;

  input                                         std__mgr51__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane13_strm1_data        ;
  output                                        mgr51__std__lane13_strm1_data_valid  ;

  input                                         std__mgr51__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane14_strm0_data        ;
  output                                        mgr51__std__lane14_strm0_data_valid  ;

  input                                         std__mgr51__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane14_strm1_data        ;
  output                                        mgr51__std__lane14_strm1_data_valid  ;

  input                                         std__mgr51__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane15_strm0_data        ;
  output                                        mgr51__std__lane15_strm0_data_valid  ;

  input                                         std__mgr51__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane15_strm1_data        ;
  output                                        mgr51__std__lane15_strm1_data_valid  ;

  input                                         std__mgr51__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane16_strm0_data        ;
  output                                        mgr51__std__lane16_strm0_data_valid  ;

  input                                         std__mgr51__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane16_strm1_data        ;
  output                                        mgr51__std__lane16_strm1_data_valid  ;

  input                                         std__mgr51__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane17_strm0_data        ;
  output                                        mgr51__std__lane17_strm0_data_valid  ;

  input                                         std__mgr51__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane17_strm1_data        ;
  output                                        mgr51__std__lane17_strm1_data_valid  ;

  input                                         std__mgr51__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane18_strm0_data        ;
  output                                        mgr51__std__lane18_strm0_data_valid  ;

  input                                         std__mgr51__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane18_strm1_data        ;
  output                                        mgr51__std__lane18_strm1_data_valid  ;

  input                                         std__mgr51__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane19_strm0_data        ;
  output                                        mgr51__std__lane19_strm0_data_valid  ;

  input                                         std__mgr51__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane19_strm1_data        ;
  output                                        mgr51__std__lane19_strm1_data_valid  ;

  input                                         std__mgr51__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane20_strm0_data        ;
  output                                        mgr51__std__lane20_strm0_data_valid  ;

  input                                         std__mgr51__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane20_strm1_data        ;
  output                                        mgr51__std__lane20_strm1_data_valid  ;

  input                                         std__mgr51__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane21_strm0_data        ;
  output                                        mgr51__std__lane21_strm0_data_valid  ;

  input                                         std__mgr51__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane21_strm1_data        ;
  output                                        mgr51__std__lane21_strm1_data_valid  ;

  input                                         std__mgr51__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane22_strm0_data        ;
  output                                        mgr51__std__lane22_strm0_data_valid  ;

  input                                         std__mgr51__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane22_strm1_data        ;
  output                                        mgr51__std__lane22_strm1_data_valid  ;

  input                                         std__mgr51__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane23_strm0_data        ;
  output                                        mgr51__std__lane23_strm0_data_valid  ;

  input                                         std__mgr51__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane23_strm1_data        ;
  output                                        mgr51__std__lane23_strm1_data_valid  ;

  input                                         std__mgr51__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane24_strm0_data        ;
  output                                        mgr51__std__lane24_strm0_data_valid  ;

  input                                         std__mgr51__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane24_strm1_data        ;
  output                                        mgr51__std__lane24_strm1_data_valid  ;

  input                                         std__mgr51__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane25_strm0_data        ;
  output                                        mgr51__std__lane25_strm0_data_valid  ;

  input                                         std__mgr51__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane25_strm1_data        ;
  output                                        mgr51__std__lane25_strm1_data_valid  ;

  input                                         std__mgr51__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane26_strm0_data        ;
  output                                        mgr51__std__lane26_strm0_data_valid  ;

  input                                         std__mgr51__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane26_strm1_data        ;
  output                                        mgr51__std__lane26_strm1_data_valid  ;

  input                                         std__mgr51__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane27_strm0_data        ;
  output                                        mgr51__std__lane27_strm0_data_valid  ;

  input                                         std__mgr51__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane27_strm1_data        ;
  output                                        mgr51__std__lane27_strm1_data_valid  ;

  input                                         std__mgr51__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane28_strm0_data        ;
  output                                        mgr51__std__lane28_strm0_data_valid  ;

  input                                         std__mgr51__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane28_strm1_data        ;
  output                                        mgr51__std__lane28_strm1_data_valid  ;

  input                                         std__mgr51__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane29_strm0_data        ;
  output                                        mgr51__std__lane29_strm0_data_valid  ;

  input                                         std__mgr51__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane29_strm1_data        ;
  output                                        mgr51__std__lane29_strm1_data_valid  ;

  input                                         std__mgr51__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane30_strm0_data        ;
  output                                        mgr51__std__lane30_strm0_data_valid  ;

  input                                         std__mgr51__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane30_strm1_data        ;
  output                                        mgr51__std__lane30_strm1_data_valid  ;

  input                                         std__mgr51__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane31_strm0_data        ;
  output                                        mgr51__std__lane31_strm0_data_valid  ;

  input                                         std__mgr51__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane31_strm1_data        ;
  output                                        mgr51__std__lane31_strm1_data_valid  ;

  input                                         std__mgr52__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane0_strm0_data        ;
  output                                        mgr52__std__lane0_strm0_data_valid  ;

  input                                         std__mgr52__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane0_strm1_data        ;
  output                                        mgr52__std__lane0_strm1_data_valid  ;

  input                                         std__mgr52__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane1_strm0_data        ;
  output                                        mgr52__std__lane1_strm0_data_valid  ;

  input                                         std__mgr52__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane1_strm1_data        ;
  output                                        mgr52__std__lane1_strm1_data_valid  ;

  input                                         std__mgr52__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane2_strm0_data        ;
  output                                        mgr52__std__lane2_strm0_data_valid  ;

  input                                         std__mgr52__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane2_strm1_data        ;
  output                                        mgr52__std__lane2_strm1_data_valid  ;

  input                                         std__mgr52__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane3_strm0_data        ;
  output                                        mgr52__std__lane3_strm0_data_valid  ;

  input                                         std__mgr52__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane3_strm1_data        ;
  output                                        mgr52__std__lane3_strm1_data_valid  ;

  input                                         std__mgr52__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane4_strm0_data        ;
  output                                        mgr52__std__lane4_strm0_data_valid  ;

  input                                         std__mgr52__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane4_strm1_data        ;
  output                                        mgr52__std__lane4_strm1_data_valid  ;

  input                                         std__mgr52__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane5_strm0_data        ;
  output                                        mgr52__std__lane5_strm0_data_valid  ;

  input                                         std__mgr52__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane5_strm1_data        ;
  output                                        mgr52__std__lane5_strm1_data_valid  ;

  input                                         std__mgr52__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane6_strm0_data        ;
  output                                        mgr52__std__lane6_strm0_data_valid  ;

  input                                         std__mgr52__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane6_strm1_data        ;
  output                                        mgr52__std__lane6_strm1_data_valid  ;

  input                                         std__mgr52__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane7_strm0_data        ;
  output                                        mgr52__std__lane7_strm0_data_valid  ;

  input                                         std__mgr52__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane7_strm1_data        ;
  output                                        mgr52__std__lane7_strm1_data_valid  ;

  input                                         std__mgr52__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane8_strm0_data        ;
  output                                        mgr52__std__lane8_strm0_data_valid  ;

  input                                         std__mgr52__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane8_strm1_data        ;
  output                                        mgr52__std__lane8_strm1_data_valid  ;

  input                                         std__mgr52__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane9_strm0_data        ;
  output                                        mgr52__std__lane9_strm0_data_valid  ;

  input                                         std__mgr52__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane9_strm1_data        ;
  output                                        mgr52__std__lane9_strm1_data_valid  ;

  input                                         std__mgr52__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane10_strm0_data        ;
  output                                        mgr52__std__lane10_strm0_data_valid  ;

  input                                         std__mgr52__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane10_strm1_data        ;
  output                                        mgr52__std__lane10_strm1_data_valid  ;

  input                                         std__mgr52__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane11_strm0_data        ;
  output                                        mgr52__std__lane11_strm0_data_valid  ;

  input                                         std__mgr52__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane11_strm1_data        ;
  output                                        mgr52__std__lane11_strm1_data_valid  ;

  input                                         std__mgr52__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane12_strm0_data        ;
  output                                        mgr52__std__lane12_strm0_data_valid  ;

  input                                         std__mgr52__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane12_strm1_data        ;
  output                                        mgr52__std__lane12_strm1_data_valid  ;

  input                                         std__mgr52__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane13_strm0_data        ;
  output                                        mgr52__std__lane13_strm0_data_valid  ;

  input                                         std__mgr52__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane13_strm1_data        ;
  output                                        mgr52__std__lane13_strm1_data_valid  ;

  input                                         std__mgr52__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane14_strm0_data        ;
  output                                        mgr52__std__lane14_strm0_data_valid  ;

  input                                         std__mgr52__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane14_strm1_data        ;
  output                                        mgr52__std__lane14_strm1_data_valid  ;

  input                                         std__mgr52__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane15_strm0_data        ;
  output                                        mgr52__std__lane15_strm0_data_valid  ;

  input                                         std__mgr52__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane15_strm1_data        ;
  output                                        mgr52__std__lane15_strm1_data_valid  ;

  input                                         std__mgr52__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane16_strm0_data        ;
  output                                        mgr52__std__lane16_strm0_data_valid  ;

  input                                         std__mgr52__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane16_strm1_data        ;
  output                                        mgr52__std__lane16_strm1_data_valid  ;

  input                                         std__mgr52__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane17_strm0_data        ;
  output                                        mgr52__std__lane17_strm0_data_valid  ;

  input                                         std__mgr52__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane17_strm1_data        ;
  output                                        mgr52__std__lane17_strm1_data_valid  ;

  input                                         std__mgr52__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane18_strm0_data        ;
  output                                        mgr52__std__lane18_strm0_data_valid  ;

  input                                         std__mgr52__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane18_strm1_data        ;
  output                                        mgr52__std__lane18_strm1_data_valid  ;

  input                                         std__mgr52__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane19_strm0_data        ;
  output                                        mgr52__std__lane19_strm0_data_valid  ;

  input                                         std__mgr52__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane19_strm1_data        ;
  output                                        mgr52__std__lane19_strm1_data_valid  ;

  input                                         std__mgr52__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane20_strm0_data        ;
  output                                        mgr52__std__lane20_strm0_data_valid  ;

  input                                         std__mgr52__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane20_strm1_data        ;
  output                                        mgr52__std__lane20_strm1_data_valid  ;

  input                                         std__mgr52__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane21_strm0_data        ;
  output                                        mgr52__std__lane21_strm0_data_valid  ;

  input                                         std__mgr52__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane21_strm1_data        ;
  output                                        mgr52__std__lane21_strm1_data_valid  ;

  input                                         std__mgr52__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane22_strm0_data        ;
  output                                        mgr52__std__lane22_strm0_data_valid  ;

  input                                         std__mgr52__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane22_strm1_data        ;
  output                                        mgr52__std__lane22_strm1_data_valid  ;

  input                                         std__mgr52__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane23_strm0_data        ;
  output                                        mgr52__std__lane23_strm0_data_valid  ;

  input                                         std__mgr52__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane23_strm1_data        ;
  output                                        mgr52__std__lane23_strm1_data_valid  ;

  input                                         std__mgr52__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane24_strm0_data        ;
  output                                        mgr52__std__lane24_strm0_data_valid  ;

  input                                         std__mgr52__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane24_strm1_data        ;
  output                                        mgr52__std__lane24_strm1_data_valid  ;

  input                                         std__mgr52__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane25_strm0_data        ;
  output                                        mgr52__std__lane25_strm0_data_valid  ;

  input                                         std__mgr52__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane25_strm1_data        ;
  output                                        mgr52__std__lane25_strm1_data_valid  ;

  input                                         std__mgr52__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane26_strm0_data        ;
  output                                        mgr52__std__lane26_strm0_data_valid  ;

  input                                         std__mgr52__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane26_strm1_data        ;
  output                                        mgr52__std__lane26_strm1_data_valid  ;

  input                                         std__mgr52__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane27_strm0_data        ;
  output                                        mgr52__std__lane27_strm0_data_valid  ;

  input                                         std__mgr52__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane27_strm1_data        ;
  output                                        mgr52__std__lane27_strm1_data_valid  ;

  input                                         std__mgr52__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane28_strm0_data        ;
  output                                        mgr52__std__lane28_strm0_data_valid  ;

  input                                         std__mgr52__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane28_strm1_data        ;
  output                                        mgr52__std__lane28_strm1_data_valid  ;

  input                                         std__mgr52__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane29_strm0_data        ;
  output                                        mgr52__std__lane29_strm0_data_valid  ;

  input                                         std__mgr52__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane29_strm1_data        ;
  output                                        mgr52__std__lane29_strm1_data_valid  ;

  input                                         std__mgr52__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane30_strm0_data        ;
  output                                        mgr52__std__lane30_strm0_data_valid  ;

  input                                         std__mgr52__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane30_strm1_data        ;
  output                                        mgr52__std__lane30_strm1_data_valid  ;

  input                                         std__mgr52__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane31_strm0_data        ;
  output                                        mgr52__std__lane31_strm0_data_valid  ;

  input                                         std__mgr52__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane31_strm1_data        ;
  output                                        mgr52__std__lane31_strm1_data_valid  ;

  input                                         std__mgr53__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane0_strm0_data        ;
  output                                        mgr53__std__lane0_strm0_data_valid  ;

  input                                         std__mgr53__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane0_strm1_data        ;
  output                                        mgr53__std__lane0_strm1_data_valid  ;

  input                                         std__mgr53__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane1_strm0_data        ;
  output                                        mgr53__std__lane1_strm0_data_valid  ;

  input                                         std__mgr53__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane1_strm1_data        ;
  output                                        mgr53__std__lane1_strm1_data_valid  ;

  input                                         std__mgr53__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane2_strm0_data        ;
  output                                        mgr53__std__lane2_strm0_data_valid  ;

  input                                         std__mgr53__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane2_strm1_data        ;
  output                                        mgr53__std__lane2_strm1_data_valid  ;

  input                                         std__mgr53__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane3_strm0_data        ;
  output                                        mgr53__std__lane3_strm0_data_valid  ;

  input                                         std__mgr53__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane3_strm1_data        ;
  output                                        mgr53__std__lane3_strm1_data_valid  ;

  input                                         std__mgr53__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane4_strm0_data        ;
  output                                        mgr53__std__lane4_strm0_data_valid  ;

  input                                         std__mgr53__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane4_strm1_data        ;
  output                                        mgr53__std__lane4_strm1_data_valid  ;

  input                                         std__mgr53__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane5_strm0_data        ;
  output                                        mgr53__std__lane5_strm0_data_valid  ;

  input                                         std__mgr53__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane5_strm1_data        ;
  output                                        mgr53__std__lane5_strm1_data_valid  ;

  input                                         std__mgr53__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane6_strm0_data        ;
  output                                        mgr53__std__lane6_strm0_data_valid  ;

  input                                         std__mgr53__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane6_strm1_data        ;
  output                                        mgr53__std__lane6_strm1_data_valid  ;

  input                                         std__mgr53__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane7_strm0_data        ;
  output                                        mgr53__std__lane7_strm0_data_valid  ;

  input                                         std__mgr53__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane7_strm1_data        ;
  output                                        mgr53__std__lane7_strm1_data_valid  ;

  input                                         std__mgr53__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane8_strm0_data        ;
  output                                        mgr53__std__lane8_strm0_data_valid  ;

  input                                         std__mgr53__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane8_strm1_data        ;
  output                                        mgr53__std__lane8_strm1_data_valid  ;

  input                                         std__mgr53__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane9_strm0_data        ;
  output                                        mgr53__std__lane9_strm0_data_valid  ;

  input                                         std__mgr53__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane9_strm1_data        ;
  output                                        mgr53__std__lane9_strm1_data_valid  ;

  input                                         std__mgr53__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane10_strm0_data        ;
  output                                        mgr53__std__lane10_strm0_data_valid  ;

  input                                         std__mgr53__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane10_strm1_data        ;
  output                                        mgr53__std__lane10_strm1_data_valid  ;

  input                                         std__mgr53__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane11_strm0_data        ;
  output                                        mgr53__std__lane11_strm0_data_valid  ;

  input                                         std__mgr53__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane11_strm1_data        ;
  output                                        mgr53__std__lane11_strm1_data_valid  ;

  input                                         std__mgr53__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane12_strm0_data        ;
  output                                        mgr53__std__lane12_strm0_data_valid  ;

  input                                         std__mgr53__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane12_strm1_data        ;
  output                                        mgr53__std__lane12_strm1_data_valid  ;

  input                                         std__mgr53__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane13_strm0_data        ;
  output                                        mgr53__std__lane13_strm0_data_valid  ;

  input                                         std__mgr53__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane13_strm1_data        ;
  output                                        mgr53__std__lane13_strm1_data_valid  ;

  input                                         std__mgr53__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane14_strm0_data        ;
  output                                        mgr53__std__lane14_strm0_data_valid  ;

  input                                         std__mgr53__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane14_strm1_data        ;
  output                                        mgr53__std__lane14_strm1_data_valid  ;

  input                                         std__mgr53__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane15_strm0_data        ;
  output                                        mgr53__std__lane15_strm0_data_valid  ;

  input                                         std__mgr53__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane15_strm1_data        ;
  output                                        mgr53__std__lane15_strm1_data_valid  ;

  input                                         std__mgr53__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane16_strm0_data        ;
  output                                        mgr53__std__lane16_strm0_data_valid  ;

  input                                         std__mgr53__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane16_strm1_data        ;
  output                                        mgr53__std__lane16_strm1_data_valid  ;

  input                                         std__mgr53__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane17_strm0_data        ;
  output                                        mgr53__std__lane17_strm0_data_valid  ;

  input                                         std__mgr53__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane17_strm1_data        ;
  output                                        mgr53__std__lane17_strm1_data_valid  ;

  input                                         std__mgr53__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane18_strm0_data        ;
  output                                        mgr53__std__lane18_strm0_data_valid  ;

  input                                         std__mgr53__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane18_strm1_data        ;
  output                                        mgr53__std__lane18_strm1_data_valid  ;

  input                                         std__mgr53__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane19_strm0_data        ;
  output                                        mgr53__std__lane19_strm0_data_valid  ;

  input                                         std__mgr53__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane19_strm1_data        ;
  output                                        mgr53__std__lane19_strm1_data_valid  ;

  input                                         std__mgr53__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane20_strm0_data        ;
  output                                        mgr53__std__lane20_strm0_data_valid  ;

  input                                         std__mgr53__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane20_strm1_data        ;
  output                                        mgr53__std__lane20_strm1_data_valid  ;

  input                                         std__mgr53__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane21_strm0_data        ;
  output                                        mgr53__std__lane21_strm0_data_valid  ;

  input                                         std__mgr53__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane21_strm1_data        ;
  output                                        mgr53__std__lane21_strm1_data_valid  ;

  input                                         std__mgr53__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane22_strm0_data        ;
  output                                        mgr53__std__lane22_strm0_data_valid  ;

  input                                         std__mgr53__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane22_strm1_data        ;
  output                                        mgr53__std__lane22_strm1_data_valid  ;

  input                                         std__mgr53__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane23_strm0_data        ;
  output                                        mgr53__std__lane23_strm0_data_valid  ;

  input                                         std__mgr53__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane23_strm1_data        ;
  output                                        mgr53__std__lane23_strm1_data_valid  ;

  input                                         std__mgr53__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane24_strm0_data        ;
  output                                        mgr53__std__lane24_strm0_data_valid  ;

  input                                         std__mgr53__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane24_strm1_data        ;
  output                                        mgr53__std__lane24_strm1_data_valid  ;

  input                                         std__mgr53__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane25_strm0_data        ;
  output                                        mgr53__std__lane25_strm0_data_valid  ;

  input                                         std__mgr53__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane25_strm1_data        ;
  output                                        mgr53__std__lane25_strm1_data_valid  ;

  input                                         std__mgr53__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane26_strm0_data        ;
  output                                        mgr53__std__lane26_strm0_data_valid  ;

  input                                         std__mgr53__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane26_strm1_data        ;
  output                                        mgr53__std__lane26_strm1_data_valid  ;

  input                                         std__mgr53__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane27_strm0_data        ;
  output                                        mgr53__std__lane27_strm0_data_valid  ;

  input                                         std__mgr53__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane27_strm1_data        ;
  output                                        mgr53__std__lane27_strm1_data_valid  ;

  input                                         std__mgr53__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane28_strm0_data        ;
  output                                        mgr53__std__lane28_strm0_data_valid  ;

  input                                         std__mgr53__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane28_strm1_data        ;
  output                                        mgr53__std__lane28_strm1_data_valid  ;

  input                                         std__mgr53__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane29_strm0_data        ;
  output                                        mgr53__std__lane29_strm0_data_valid  ;

  input                                         std__mgr53__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane29_strm1_data        ;
  output                                        mgr53__std__lane29_strm1_data_valid  ;

  input                                         std__mgr53__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane30_strm0_data        ;
  output                                        mgr53__std__lane30_strm0_data_valid  ;

  input                                         std__mgr53__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane30_strm1_data        ;
  output                                        mgr53__std__lane30_strm1_data_valid  ;

  input                                         std__mgr53__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane31_strm0_data        ;
  output                                        mgr53__std__lane31_strm0_data_valid  ;

  input                                         std__mgr53__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane31_strm1_data        ;
  output                                        mgr53__std__lane31_strm1_data_valid  ;

  input                                         std__mgr54__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane0_strm0_data        ;
  output                                        mgr54__std__lane0_strm0_data_valid  ;

  input                                         std__mgr54__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane0_strm1_data        ;
  output                                        mgr54__std__lane0_strm1_data_valid  ;

  input                                         std__mgr54__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane1_strm0_data        ;
  output                                        mgr54__std__lane1_strm0_data_valid  ;

  input                                         std__mgr54__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane1_strm1_data        ;
  output                                        mgr54__std__lane1_strm1_data_valid  ;

  input                                         std__mgr54__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane2_strm0_data        ;
  output                                        mgr54__std__lane2_strm0_data_valid  ;

  input                                         std__mgr54__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane2_strm1_data        ;
  output                                        mgr54__std__lane2_strm1_data_valid  ;

  input                                         std__mgr54__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane3_strm0_data        ;
  output                                        mgr54__std__lane3_strm0_data_valid  ;

  input                                         std__mgr54__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane3_strm1_data        ;
  output                                        mgr54__std__lane3_strm1_data_valid  ;

  input                                         std__mgr54__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane4_strm0_data        ;
  output                                        mgr54__std__lane4_strm0_data_valid  ;

  input                                         std__mgr54__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane4_strm1_data        ;
  output                                        mgr54__std__lane4_strm1_data_valid  ;

  input                                         std__mgr54__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane5_strm0_data        ;
  output                                        mgr54__std__lane5_strm0_data_valid  ;

  input                                         std__mgr54__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane5_strm1_data        ;
  output                                        mgr54__std__lane5_strm1_data_valid  ;

  input                                         std__mgr54__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane6_strm0_data        ;
  output                                        mgr54__std__lane6_strm0_data_valid  ;

  input                                         std__mgr54__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane6_strm1_data        ;
  output                                        mgr54__std__lane6_strm1_data_valid  ;

  input                                         std__mgr54__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane7_strm0_data        ;
  output                                        mgr54__std__lane7_strm0_data_valid  ;

  input                                         std__mgr54__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane7_strm1_data        ;
  output                                        mgr54__std__lane7_strm1_data_valid  ;

  input                                         std__mgr54__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane8_strm0_data        ;
  output                                        mgr54__std__lane8_strm0_data_valid  ;

  input                                         std__mgr54__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane8_strm1_data        ;
  output                                        mgr54__std__lane8_strm1_data_valid  ;

  input                                         std__mgr54__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane9_strm0_data        ;
  output                                        mgr54__std__lane9_strm0_data_valid  ;

  input                                         std__mgr54__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane9_strm1_data        ;
  output                                        mgr54__std__lane9_strm1_data_valid  ;

  input                                         std__mgr54__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane10_strm0_data        ;
  output                                        mgr54__std__lane10_strm0_data_valid  ;

  input                                         std__mgr54__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane10_strm1_data        ;
  output                                        mgr54__std__lane10_strm1_data_valid  ;

  input                                         std__mgr54__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane11_strm0_data        ;
  output                                        mgr54__std__lane11_strm0_data_valid  ;

  input                                         std__mgr54__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane11_strm1_data        ;
  output                                        mgr54__std__lane11_strm1_data_valid  ;

  input                                         std__mgr54__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane12_strm0_data        ;
  output                                        mgr54__std__lane12_strm0_data_valid  ;

  input                                         std__mgr54__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane12_strm1_data        ;
  output                                        mgr54__std__lane12_strm1_data_valid  ;

  input                                         std__mgr54__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane13_strm0_data        ;
  output                                        mgr54__std__lane13_strm0_data_valid  ;

  input                                         std__mgr54__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane13_strm1_data        ;
  output                                        mgr54__std__lane13_strm1_data_valid  ;

  input                                         std__mgr54__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane14_strm0_data        ;
  output                                        mgr54__std__lane14_strm0_data_valid  ;

  input                                         std__mgr54__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane14_strm1_data        ;
  output                                        mgr54__std__lane14_strm1_data_valid  ;

  input                                         std__mgr54__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane15_strm0_data        ;
  output                                        mgr54__std__lane15_strm0_data_valid  ;

  input                                         std__mgr54__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane15_strm1_data        ;
  output                                        mgr54__std__lane15_strm1_data_valid  ;

  input                                         std__mgr54__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane16_strm0_data        ;
  output                                        mgr54__std__lane16_strm0_data_valid  ;

  input                                         std__mgr54__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane16_strm1_data        ;
  output                                        mgr54__std__lane16_strm1_data_valid  ;

  input                                         std__mgr54__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane17_strm0_data        ;
  output                                        mgr54__std__lane17_strm0_data_valid  ;

  input                                         std__mgr54__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane17_strm1_data        ;
  output                                        mgr54__std__lane17_strm1_data_valid  ;

  input                                         std__mgr54__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane18_strm0_data        ;
  output                                        mgr54__std__lane18_strm0_data_valid  ;

  input                                         std__mgr54__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane18_strm1_data        ;
  output                                        mgr54__std__lane18_strm1_data_valid  ;

  input                                         std__mgr54__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane19_strm0_data        ;
  output                                        mgr54__std__lane19_strm0_data_valid  ;

  input                                         std__mgr54__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane19_strm1_data        ;
  output                                        mgr54__std__lane19_strm1_data_valid  ;

  input                                         std__mgr54__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane20_strm0_data        ;
  output                                        mgr54__std__lane20_strm0_data_valid  ;

  input                                         std__mgr54__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane20_strm1_data        ;
  output                                        mgr54__std__lane20_strm1_data_valid  ;

  input                                         std__mgr54__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane21_strm0_data        ;
  output                                        mgr54__std__lane21_strm0_data_valid  ;

  input                                         std__mgr54__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane21_strm1_data        ;
  output                                        mgr54__std__lane21_strm1_data_valid  ;

  input                                         std__mgr54__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane22_strm0_data        ;
  output                                        mgr54__std__lane22_strm0_data_valid  ;

  input                                         std__mgr54__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane22_strm1_data        ;
  output                                        mgr54__std__lane22_strm1_data_valid  ;

  input                                         std__mgr54__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane23_strm0_data        ;
  output                                        mgr54__std__lane23_strm0_data_valid  ;

  input                                         std__mgr54__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane23_strm1_data        ;
  output                                        mgr54__std__lane23_strm1_data_valid  ;

  input                                         std__mgr54__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane24_strm0_data        ;
  output                                        mgr54__std__lane24_strm0_data_valid  ;

  input                                         std__mgr54__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane24_strm1_data        ;
  output                                        mgr54__std__lane24_strm1_data_valid  ;

  input                                         std__mgr54__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane25_strm0_data        ;
  output                                        mgr54__std__lane25_strm0_data_valid  ;

  input                                         std__mgr54__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane25_strm1_data        ;
  output                                        mgr54__std__lane25_strm1_data_valid  ;

  input                                         std__mgr54__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane26_strm0_data        ;
  output                                        mgr54__std__lane26_strm0_data_valid  ;

  input                                         std__mgr54__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane26_strm1_data        ;
  output                                        mgr54__std__lane26_strm1_data_valid  ;

  input                                         std__mgr54__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane27_strm0_data        ;
  output                                        mgr54__std__lane27_strm0_data_valid  ;

  input                                         std__mgr54__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane27_strm1_data        ;
  output                                        mgr54__std__lane27_strm1_data_valid  ;

  input                                         std__mgr54__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane28_strm0_data        ;
  output                                        mgr54__std__lane28_strm0_data_valid  ;

  input                                         std__mgr54__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane28_strm1_data        ;
  output                                        mgr54__std__lane28_strm1_data_valid  ;

  input                                         std__mgr54__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane29_strm0_data        ;
  output                                        mgr54__std__lane29_strm0_data_valid  ;

  input                                         std__mgr54__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane29_strm1_data        ;
  output                                        mgr54__std__lane29_strm1_data_valid  ;

  input                                         std__mgr54__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane30_strm0_data        ;
  output                                        mgr54__std__lane30_strm0_data_valid  ;

  input                                         std__mgr54__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane30_strm1_data        ;
  output                                        mgr54__std__lane30_strm1_data_valid  ;

  input                                         std__mgr54__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane31_strm0_data        ;
  output                                        mgr54__std__lane31_strm0_data_valid  ;

  input                                         std__mgr54__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane31_strm1_data        ;
  output                                        mgr54__std__lane31_strm1_data_valid  ;

  input                                         std__mgr55__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane0_strm0_data        ;
  output                                        mgr55__std__lane0_strm0_data_valid  ;

  input                                         std__mgr55__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane0_strm1_data        ;
  output                                        mgr55__std__lane0_strm1_data_valid  ;

  input                                         std__mgr55__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane1_strm0_data        ;
  output                                        mgr55__std__lane1_strm0_data_valid  ;

  input                                         std__mgr55__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane1_strm1_data        ;
  output                                        mgr55__std__lane1_strm1_data_valid  ;

  input                                         std__mgr55__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane2_strm0_data        ;
  output                                        mgr55__std__lane2_strm0_data_valid  ;

  input                                         std__mgr55__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane2_strm1_data        ;
  output                                        mgr55__std__lane2_strm1_data_valid  ;

  input                                         std__mgr55__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane3_strm0_data        ;
  output                                        mgr55__std__lane3_strm0_data_valid  ;

  input                                         std__mgr55__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane3_strm1_data        ;
  output                                        mgr55__std__lane3_strm1_data_valid  ;

  input                                         std__mgr55__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane4_strm0_data        ;
  output                                        mgr55__std__lane4_strm0_data_valid  ;

  input                                         std__mgr55__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane4_strm1_data        ;
  output                                        mgr55__std__lane4_strm1_data_valid  ;

  input                                         std__mgr55__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane5_strm0_data        ;
  output                                        mgr55__std__lane5_strm0_data_valid  ;

  input                                         std__mgr55__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane5_strm1_data        ;
  output                                        mgr55__std__lane5_strm1_data_valid  ;

  input                                         std__mgr55__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane6_strm0_data        ;
  output                                        mgr55__std__lane6_strm0_data_valid  ;

  input                                         std__mgr55__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane6_strm1_data        ;
  output                                        mgr55__std__lane6_strm1_data_valid  ;

  input                                         std__mgr55__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane7_strm0_data        ;
  output                                        mgr55__std__lane7_strm0_data_valid  ;

  input                                         std__mgr55__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane7_strm1_data        ;
  output                                        mgr55__std__lane7_strm1_data_valid  ;

  input                                         std__mgr55__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane8_strm0_data        ;
  output                                        mgr55__std__lane8_strm0_data_valid  ;

  input                                         std__mgr55__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane8_strm1_data        ;
  output                                        mgr55__std__lane8_strm1_data_valid  ;

  input                                         std__mgr55__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane9_strm0_data        ;
  output                                        mgr55__std__lane9_strm0_data_valid  ;

  input                                         std__mgr55__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane9_strm1_data        ;
  output                                        mgr55__std__lane9_strm1_data_valid  ;

  input                                         std__mgr55__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane10_strm0_data        ;
  output                                        mgr55__std__lane10_strm0_data_valid  ;

  input                                         std__mgr55__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane10_strm1_data        ;
  output                                        mgr55__std__lane10_strm1_data_valid  ;

  input                                         std__mgr55__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane11_strm0_data        ;
  output                                        mgr55__std__lane11_strm0_data_valid  ;

  input                                         std__mgr55__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane11_strm1_data        ;
  output                                        mgr55__std__lane11_strm1_data_valid  ;

  input                                         std__mgr55__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane12_strm0_data        ;
  output                                        mgr55__std__lane12_strm0_data_valid  ;

  input                                         std__mgr55__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane12_strm1_data        ;
  output                                        mgr55__std__lane12_strm1_data_valid  ;

  input                                         std__mgr55__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane13_strm0_data        ;
  output                                        mgr55__std__lane13_strm0_data_valid  ;

  input                                         std__mgr55__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane13_strm1_data        ;
  output                                        mgr55__std__lane13_strm1_data_valid  ;

  input                                         std__mgr55__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane14_strm0_data        ;
  output                                        mgr55__std__lane14_strm0_data_valid  ;

  input                                         std__mgr55__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane14_strm1_data        ;
  output                                        mgr55__std__lane14_strm1_data_valid  ;

  input                                         std__mgr55__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane15_strm0_data        ;
  output                                        mgr55__std__lane15_strm0_data_valid  ;

  input                                         std__mgr55__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane15_strm1_data        ;
  output                                        mgr55__std__lane15_strm1_data_valid  ;

  input                                         std__mgr55__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane16_strm0_data        ;
  output                                        mgr55__std__lane16_strm0_data_valid  ;

  input                                         std__mgr55__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane16_strm1_data        ;
  output                                        mgr55__std__lane16_strm1_data_valid  ;

  input                                         std__mgr55__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane17_strm0_data        ;
  output                                        mgr55__std__lane17_strm0_data_valid  ;

  input                                         std__mgr55__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane17_strm1_data        ;
  output                                        mgr55__std__lane17_strm1_data_valid  ;

  input                                         std__mgr55__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane18_strm0_data        ;
  output                                        mgr55__std__lane18_strm0_data_valid  ;

  input                                         std__mgr55__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane18_strm1_data        ;
  output                                        mgr55__std__lane18_strm1_data_valid  ;

  input                                         std__mgr55__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane19_strm0_data        ;
  output                                        mgr55__std__lane19_strm0_data_valid  ;

  input                                         std__mgr55__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane19_strm1_data        ;
  output                                        mgr55__std__lane19_strm1_data_valid  ;

  input                                         std__mgr55__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane20_strm0_data        ;
  output                                        mgr55__std__lane20_strm0_data_valid  ;

  input                                         std__mgr55__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane20_strm1_data        ;
  output                                        mgr55__std__lane20_strm1_data_valid  ;

  input                                         std__mgr55__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane21_strm0_data        ;
  output                                        mgr55__std__lane21_strm0_data_valid  ;

  input                                         std__mgr55__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane21_strm1_data        ;
  output                                        mgr55__std__lane21_strm1_data_valid  ;

  input                                         std__mgr55__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane22_strm0_data        ;
  output                                        mgr55__std__lane22_strm0_data_valid  ;

  input                                         std__mgr55__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane22_strm1_data        ;
  output                                        mgr55__std__lane22_strm1_data_valid  ;

  input                                         std__mgr55__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane23_strm0_data        ;
  output                                        mgr55__std__lane23_strm0_data_valid  ;

  input                                         std__mgr55__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane23_strm1_data        ;
  output                                        mgr55__std__lane23_strm1_data_valid  ;

  input                                         std__mgr55__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane24_strm0_data        ;
  output                                        mgr55__std__lane24_strm0_data_valid  ;

  input                                         std__mgr55__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane24_strm1_data        ;
  output                                        mgr55__std__lane24_strm1_data_valid  ;

  input                                         std__mgr55__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane25_strm0_data        ;
  output                                        mgr55__std__lane25_strm0_data_valid  ;

  input                                         std__mgr55__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane25_strm1_data        ;
  output                                        mgr55__std__lane25_strm1_data_valid  ;

  input                                         std__mgr55__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane26_strm0_data        ;
  output                                        mgr55__std__lane26_strm0_data_valid  ;

  input                                         std__mgr55__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane26_strm1_data        ;
  output                                        mgr55__std__lane26_strm1_data_valid  ;

  input                                         std__mgr55__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane27_strm0_data        ;
  output                                        mgr55__std__lane27_strm0_data_valid  ;

  input                                         std__mgr55__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane27_strm1_data        ;
  output                                        mgr55__std__lane27_strm1_data_valid  ;

  input                                         std__mgr55__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane28_strm0_data        ;
  output                                        mgr55__std__lane28_strm0_data_valid  ;

  input                                         std__mgr55__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane28_strm1_data        ;
  output                                        mgr55__std__lane28_strm1_data_valid  ;

  input                                         std__mgr55__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane29_strm0_data        ;
  output                                        mgr55__std__lane29_strm0_data_valid  ;

  input                                         std__mgr55__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane29_strm1_data        ;
  output                                        mgr55__std__lane29_strm1_data_valid  ;

  input                                         std__mgr55__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane30_strm0_data        ;
  output                                        mgr55__std__lane30_strm0_data_valid  ;

  input                                         std__mgr55__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane30_strm1_data        ;
  output                                        mgr55__std__lane30_strm1_data_valid  ;

  input                                         std__mgr55__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane31_strm0_data        ;
  output                                        mgr55__std__lane31_strm0_data_valid  ;

  input                                         std__mgr55__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane31_strm1_data        ;
  output                                        mgr55__std__lane31_strm1_data_valid  ;

  input                                         std__mgr56__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane0_strm0_data        ;
  output                                        mgr56__std__lane0_strm0_data_valid  ;

  input                                         std__mgr56__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane0_strm1_data        ;
  output                                        mgr56__std__lane0_strm1_data_valid  ;

  input                                         std__mgr56__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane1_strm0_data        ;
  output                                        mgr56__std__lane1_strm0_data_valid  ;

  input                                         std__mgr56__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane1_strm1_data        ;
  output                                        mgr56__std__lane1_strm1_data_valid  ;

  input                                         std__mgr56__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane2_strm0_data        ;
  output                                        mgr56__std__lane2_strm0_data_valid  ;

  input                                         std__mgr56__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane2_strm1_data        ;
  output                                        mgr56__std__lane2_strm1_data_valid  ;

  input                                         std__mgr56__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane3_strm0_data        ;
  output                                        mgr56__std__lane3_strm0_data_valid  ;

  input                                         std__mgr56__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane3_strm1_data        ;
  output                                        mgr56__std__lane3_strm1_data_valid  ;

  input                                         std__mgr56__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane4_strm0_data        ;
  output                                        mgr56__std__lane4_strm0_data_valid  ;

  input                                         std__mgr56__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane4_strm1_data        ;
  output                                        mgr56__std__lane4_strm1_data_valid  ;

  input                                         std__mgr56__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane5_strm0_data        ;
  output                                        mgr56__std__lane5_strm0_data_valid  ;

  input                                         std__mgr56__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane5_strm1_data        ;
  output                                        mgr56__std__lane5_strm1_data_valid  ;

  input                                         std__mgr56__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane6_strm0_data        ;
  output                                        mgr56__std__lane6_strm0_data_valid  ;

  input                                         std__mgr56__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane6_strm1_data        ;
  output                                        mgr56__std__lane6_strm1_data_valid  ;

  input                                         std__mgr56__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane7_strm0_data        ;
  output                                        mgr56__std__lane7_strm0_data_valid  ;

  input                                         std__mgr56__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane7_strm1_data        ;
  output                                        mgr56__std__lane7_strm1_data_valid  ;

  input                                         std__mgr56__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane8_strm0_data        ;
  output                                        mgr56__std__lane8_strm0_data_valid  ;

  input                                         std__mgr56__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane8_strm1_data        ;
  output                                        mgr56__std__lane8_strm1_data_valid  ;

  input                                         std__mgr56__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane9_strm0_data        ;
  output                                        mgr56__std__lane9_strm0_data_valid  ;

  input                                         std__mgr56__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane9_strm1_data        ;
  output                                        mgr56__std__lane9_strm1_data_valid  ;

  input                                         std__mgr56__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane10_strm0_data        ;
  output                                        mgr56__std__lane10_strm0_data_valid  ;

  input                                         std__mgr56__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane10_strm1_data        ;
  output                                        mgr56__std__lane10_strm1_data_valid  ;

  input                                         std__mgr56__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane11_strm0_data        ;
  output                                        mgr56__std__lane11_strm0_data_valid  ;

  input                                         std__mgr56__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane11_strm1_data        ;
  output                                        mgr56__std__lane11_strm1_data_valid  ;

  input                                         std__mgr56__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane12_strm0_data        ;
  output                                        mgr56__std__lane12_strm0_data_valid  ;

  input                                         std__mgr56__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane12_strm1_data        ;
  output                                        mgr56__std__lane12_strm1_data_valid  ;

  input                                         std__mgr56__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane13_strm0_data        ;
  output                                        mgr56__std__lane13_strm0_data_valid  ;

  input                                         std__mgr56__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane13_strm1_data        ;
  output                                        mgr56__std__lane13_strm1_data_valid  ;

  input                                         std__mgr56__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane14_strm0_data        ;
  output                                        mgr56__std__lane14_strm0_data_valid  ;

  input                                         std__mgr56__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane14_strm1_data        ;
  output                                        mgr56__std__lane14_strm1_data_valid  ;

  input                                         std__mgr56__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane15_strm0_data        ;
  output                                        mgr56__std__lane15_strm0_data_valid  ;

  input                                         std__mgr56__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane15_strm1_data        ;
  output                                        mgr56__std__lane15_strm1_data_valid  ;

  input                                         std__mgr56__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane16_strm0_data        ;
  output                                        mgr56__std__lane16_strm0_data_valid  ;

  input                                         std__mgr56__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane16_strm1_data        ;
  output                                        mgr56__std__lane16_strm1_data_valid  ;

  input                                         std__mgr56__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane17_strm0_data        ;
  output                                        mgr56__std__lane17_strm0_data_valid  ;

  input                                         std__mgr56__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane17_strm1_data        ;
  output                                        mgr56__std__lane17_strm1_data_valid  ;

  input                                         std__mgr56__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane18_strm0_data        ;
  output                                        mgr56__std__lane18_strm0_data_valid  ;

  input                                         std__mgr56__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane18_strm1_data        ;
  output                                        mgr56__std__lane18_strm1_data_valid  ;

  input                                         std__mgr56__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane19_strm0_data        ;
  output                                        mgr56__std__lane19_strm0_data_valid  ;

  input                                         std__mgr56__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane19_strm1_data        ;
  output                                        mgr56__std__lane19_strm1_data_valid  ;

  input                                         std__mgr56__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane20_strm0_data        ;
  output                                        mgr56__std__lane20_strm0_data_valid  ;

  input                                         std__mgr56__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane20_strm1_data        ;
  output                                        mgr56__std__lane20_strm1_data_valid  ;

  input                                         std__mgr56__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane21_strm0_data        ;
  output                                        mgr56__std__lane21_strm0_data_valid  ;

  input                                         std__mgr56__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane21_strm1_data        ;
  output                                        mgr56__std__lane21_strm1_data_valid  ;

  input                                         std__mgr56__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane22_strm0_data        ;
  output                                        mgr56__std__lane22_strm0_data_valid  ;

  input                                         std__mgr56__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane22_strm1_data        ;
  output                                        mgr56__std__lane22_strm1_data_valid  ;

  input                                         std__mgr56__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane23_strm0_data        ;
  output                                        mgr56__std__lane23_strm0_data_valid  ;

  input                                         std__mgr56__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane23_strm1_data        ;
  output                                        mgr56__std__lane23_strm1_data_valid  ;

  input                                         std__mgr56__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane24_strm0_data        ;
  output                                        mgr56__std__lane24_strm0_data_valid  ;

  input                                         std__mgr56__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane24_strm1_data        ;
  output                                        mgr56__std__lane24_strm1_data_valid  ;

  input                                         std__mgr56__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane25_strm0_data        ;
  output                                        mgr56__std__lane25_strm0_data_valid  ;

  input                                         std__mgr56__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane25_strm1_data        ;
  output                                        mgr56__std__lane25_strm1_data_valid  ;

  input                                         std__mgr56__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane26_strm0_data        ;
  output                                        mgr56__std__lane26_strm0_data_valid  ;

  input                                         std__mgr56__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane26_strm1_data        ;
  output                                        mgr56__std__lane26_strm1_data_valid  ;

  input                                         std__mgr56__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane27_strm0_data        ;
  output                                        mgr56__std__lane27_strm0_data_valid  ;

  input                                         std__mgr56__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane27_strm1_data        ;
  output                                        mgr56__std__lane27_strm1_data_valid  ;

  input                                         std__mgr56__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane28_strm0_data        ;
  output                                        mgr56__std__lane28_strm0_data_valid  ;

  input                                         std__mgr56__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane28_strm1_data        ;
  output                                        mgr56__std__lane28_strm1_data_valid  ;

  input                                         std__mgr56__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane29_strm0_data        ;
  output                                        mgr56__std__lane29_strm0_data_valid  ;

  input                                         std__mgr56__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane29_strm1_data        ;
  output                                        mgr56__std__lane29_strm1_data_valid  ;

  input                                         std__mgr56__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane30_strm0_data        ;
  output                                        mgr56__std__lane30_strm0_data_valid  ;

  input                                         std__mgr56__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane30_strm1_data        ;
  output                                        mgr56__std__lane30_strm1_data_valid  ;

  input                                         std__mgr56__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane31_strm0_data        ;
  output                                        mgr56__std__lane31_strm0_data_valid  ;

  input                                         std__mgr56__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane31_strm1_data        ;
  output                                        mgr56__std__lane31_strm1_data_valid  ;

  input                                         std__mgr57__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane0_strm0_data        ;
  output                                        mgr57__std__lane0_strm0_data_valid  ;

  input                                         std__mgr57__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane0_strm1_data        ;
  output                                        mgr57__std__lane0_strm1_data_valid  ;

  input                                         std__mgr57__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane1_strm0_data        ;
  output                                        mgr57__std__lane1_strm0_data_valid  ;

  input                                         std__mgr57__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane1_strm1_data        ;
  output                                        mgr57__std__lane1_strm1_data_valid  ;

  input                                         std__mgr57__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane2_strm0_data        ;
  output                                        mgr57__std__lane2_strm0_data_valid  ;

  input                                         std__mgr57__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane2_strm1_data        ;
  output                                        mgr57__std__lane2_strm1_data_valid  ;

  input                                         std__mgr57__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane3_strm0_data        ;
  output                                        mgr57__std__lane3_strm0_data_valid  ;

  input                                         std__mgr57__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane3_strm1_data        ;
  output                                        mgr57__std__lane3_strm1_data_valid  ;

  input                                         std__mgr57__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane4_strm0_data        ;
  output                                        mgr57__std__lane4_strm0_data_valid  ;

  input                                         std__mgr57__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane4_strm1_data        ;
  output                                        mgr57__std__lane4_strm1_data_valid  ;

  input                                         std__mgr57__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane5_strm0_data        ;
  output                                        mgr57__std__lane5_strm0_data_valid  ;

  input                                         std__mgr57__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane5_strm1_data        ;
  output                                        mgr57__std__lane5_strm1_data_valid  ;

  input                                         std__mgr57__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane6_strm0_data        ;
  output                                        mgr57__std__lane6_strm0_data_valid  ;

  input                                         std__mgr57__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane6_strm1_data        ;
  output                                        mgr57__std__lane6_strm1_data_valid  ;

  input                                         std__mgr57__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane7_strm0_data        ;
  output                                        mgr57__std__lane7_strm0_data_valid  ;

  input                                         std__mgr57__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane7_strm1_data        ;
  output                                        mgr57__std__lane7_strm1_data_valid  ;

  input                                         std__mgr57__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane8_strm0_data        ;
  output                                        mgr57__std__lane8_strm0_data_valid  ;

  input                                         std__mgr57__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane8_strm1_data        ;
  output                                        mgr57__std__lane8_strm1_data_valid  ;

  input                                         std__mgr57__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane9_strm0_data        ;
  output                                        mgr57__std__lane9_strm0_data_valid  ;

  input                                         std__mgr57__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane9_strm1_data        ;
  output                                        mgr57__std__lane9_strm1_data_valid  ;

  input                                         std__mgr57__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane10_strm0_data        ;
  output                                        mgr57__std__lane10_strm0_data_valid  ;

  input                                         std__mgr57__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane10_strm1_data        ;
  output                                        mgr57__std__lane10_strm1_data_valid  ;

  input                                         std__mgr57__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane11_strm0_data        ;
  output                                        mgr57__std__lane11_strm0_data_valid  ;

  input                                         std__mgr57__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane11_strm1_data        ;
  output                                        mgr57__std__lane11_strm1_data_valid  ;

  input                                         std__mgr57__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane12_strm0_data        ;
  output                                        mgr57__std__lane12_strm0_data_valid  ;

  input                                         std__mgr57__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane12_strm1_data        ;
  output                                        mgr57__std__lane12_strm1_data_valid  ;

  input                                         std__mgr57__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane13_strm0_data        ;
  output                                        mgr57__std__lane13_strm0_data_valid  ;

  input                                         std__mgr57__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane13_strm1_data        ;
  output                                        mgr57__std__lane13_strm1_data_valid  ;

  input                                         std__mgr57__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane14_strm0_data        ;
  output                                        mgr57__std__lane14_strm0_data_valid  ;

  input                                         std__mgr57__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane14_strm1_data        ;
  output                                        mgr57__std__lane14_strm1_data_valid  ;

  input                                         std__mgr57__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane15_strm0_data        ;
  output                                        mgr57__std__lane15_strm0_data_valid  ;

  input                                         std__mgr57__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane15_strm1_data        ;
  output                                        mgr57__std__lane15_strm1_data_valid  ;

  input                                         std__mgr57__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane16_strm0_data        ;
  output                                        mgr57__std__lane16_strm0_data_valid  ;

  input                                         std__mgr57__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane16_strm1_data        ;
  output                                        mgr57__std__lane16_strm1_data_valid  ;

  input                                         std__mgr57__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane17_strm0_data        ;
  output                                        mgr57__std__lane17_strm0_data_valid  ;

  input                                         std__mgr57__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane17_strm1_data        ;
  output                                        mgr57__std__lane17_strm1_data_valid  ;

  input                                         std__mgr57__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane18_strm0_data        ;
  output                                        mgr57__std__lane18_strm0_data_valid  ;

  input                                         std__mgr57__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane18_strm1_data        ;
  output                                        mgr57__std__lane18_strm1_data_valid  ;

  input                                         std__mgr57__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane19_strm0_data        ;
  output                                        mgr57__std__lane19_strm0_data_valid  ;

  input                                         std__mgr57__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane19_strm1_data        ;
  output                                        mgr57__std__lane19_strm1_data_valid  ;

  input                                         std__mgr57__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane20_strm0_data        ;
  output                                        mgr57__std__lane20_strm0_data_valid  ;

  input                                         std__mgr57__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane20_strm1_data        ;
  output                                        mgr57__std__lane20_strm1_data_valid  ;

  input                                         std__mgr57__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane21_strm0_data        ;
  output                                        mgr57__std__lane21_strm0_data_valid  ;

  input                                         std__mgr57__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane21_strm1_data        ;
  output                                        mgr57__std__lane21_strm1_data_valid  ;

  input                                         std__mgr57__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane22_strm0_data        ;
  output                                        mgr57__std__lane22_strm0_data_valid  ;

  input                                         std__mgr57__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane22_strm1_data        ;
  output                                        mgr57__std__lane22_strm1_data_valid  ;

  input                                         std__mgr57__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane23_strm0_data        ;
  output                                        mgr57__std__lane23_strm0_data_valid  ;

  input                                         std__mgr57__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane23_strm1_data        ;
  output                                        mgr57__std__lane23_strm1_data_valid  ;

  input                                         std__mgr57__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane24_strm0_data        ;
  output                                        mgr57__std__lane24_strm0_data_valid  ;

  input                                         std__mgr57__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane24_strm1_data        ;
  output                                        mgr57__std__lane24_strm1_data_valid  ;

  input                                         std__mgr57__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane25_strm0_data        ;
  output                                        mgr57__std__lane25_strm0_data_valid  ;

  input                                         std__mgr57__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane25_strm1_data        ;
  output                                        mgr57__std__lane25_strm1_data_valid  ;

  input                                         std__mgr57__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane26_strm0_data        ;
  output                                        mgr57__std__lane26_strm0_data_valid  ;

  input                                         std__mgr57__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane26_strm1_data        ;
  output                                        mgr57__std__lane26_strm1_data_valid  ;

  input                                         std__mgr57__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane27_strm0_data        ;
  output                                        mgr57__std__lane27_strm0_data_valid  ;

  input                                         std__mgr57__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane27_strm1_data        ;
  output                                        mgr57__std__lane27_strm1_data_valid  ;

  input                                         std__mgr57__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane28_strm0_data        ;
  output                                        mgr57__std__lane28_strm0_data_valid  ;

  input                                         std__mgr57__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane28_strm1_data        ;
  output                                        mgr57__std__lane28_strm1_data_valid  ;

  input                                         std__mgr57__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane29_strm0_data        ;
  output                                        mgr57__std__lane29_strm0_data_valid  ;

  input                                         std__mgr57__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane29_strm1_data        ;
  output                                        mgr57__std__lane29_strm1_data_valid  ;

  input                                         std__mgr57__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane30_strm0_data        ;
  output                                        mgr57__std__lane30_strm0_data_valid  ;

  input                                         std__mgr57__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane30_strm1_data        ;
  output                                        mgr57__std__lane30_strm1_data_valid  ;

  input                                         std__mgr57__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane31_strm0_data        ;
  output                                        mgr57__std__lane31_strm0_data_valid  ;

  input                                         std__mgr57__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane31_strm1_data        ;
  output                                        mgr57__std__lane31_strm1_data_valid  ;

  input                                         std__mgr58__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane0_strm0_data        ;
  output                                        mgr58__std__lane0_strm0_data_valid  ;

  input                                         std__mgr58__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane0_strm1_data        ;
  output                                        mgr58__std__lane0_strm1_data_valid  ;

  input                                         std__mgr58__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane1_strm0_data        ;
  output                                        mgr58__std__lane1_strm0_data_valid  ;

  input                                         std__mgr58__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane1_strm1_data        ;
  output                                        mgr58__std__lane1_strm1_data_valid  ;

  input                                         std__mgr58__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane2_strm0_data        ;
  output                                        mgr58__std__lane2_strm0_data_valid  ;

  input                                         std__mgr58__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane2_strm1_data        ;
  output                                        mgr58__std__lane2_strm1_data_valid  ;

  input                                         std__mgr58__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane3_strm0_data        ;
  output                                        mgr58__std__lane3_strm0_data_valid  ;

  input                                         std__mgr58__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane3_strm1_data        ;
  output                                        mgr58__std__lane3_strm1_data_valid  ;

  input                                         std__mgr58__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane4_strm0_data        ;
  output                                        mgr58__std__lane4_strm0_data_valid  ;

  input                                         std__mgr58__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane4_strm1_data        ;
  output                                        mgr58__std__lane4_strm1_data_valid  ;

  input                                         std__mgr58__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane5_strm0_data        ;
  output                                        mgr58__std__lane5_strm0_data_valid  ;

  input                                         std__mgr58__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane5_strm1_data        ;
  output                                        mgr58__std__lane5_strm1_data_valid  ;

  input                                         std__mgr58__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane6_strm0_data        ;
  output                                        mgr58__std__lane6_strm0_data_valid  ;

  input                                         std__mgr58__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane6_strm1_data        ;
  output                                        mgr58__std__lane6_strm1_data_valid  ;

  input                                         std__mgr58__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane7_strm0_data        ;
  output                                        mgr58__std__lane7_strm0_data_valid  ;

  input                                         std__mgr58__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane7_strm1_data        ;
  output                                        mgr58__std__lane7_strm1_data_valid  ;

  input                                         std__mgr58__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane8_strm0_data        ;
  output                                        mgr58__std__lane8_strm0_data_valid  ;

  input                                         std__mgr58__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane8_strm1_data        ;
  output                                        mgr58__std__lane8_strm1_data_valid  ;

  input                                         std__mgr58__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane9_strm0_data        ;
  output                                        mgr58__std__lane9_strm0_data_valid  ;

  input                                         std__mgr58__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane9_strm1_data        ;
  output                                        mgr58__std__lane9_strm1_data_valid  ;

  input                                         std__mgr58__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane10_strm0_data        ;
  output                                        mgr58__std__lane10_strm0_data_valid  ;

  input                                         std__mgr58__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane10_strm1_data        ;
  output                                        mgr58__std__lane10_strm1_data_valid  ;

  input                                         std__mgr58__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane11_strm0_data        ;
  output                                        mgr58__std__lane11_strm0_data_valid  ;

  input                                         std__mgr58__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane11_strm1_data        ;
  output                                        mgr58__std__lane11_strm1_data_valid  ;

  input                                         std__mgr58__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane12_strm0_data        ;
  output                                        mgr58__std__lane12_strm0_data_valid  ;

  input                                         std__mgr58__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane12_strm1_data        ;
  output                                        mgr58__std__lane12_strm1_data_valid  ;

  input                                         std__mgr58__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane13_strm0_data        ;
  output                                        mgr58__std__lane13_strm0_data_valid  ;

  input                                         std__mgr58__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane13_strm1_data        ;
  output                                        mgr58__std__lane13_strm1_data_valid  ;

  input                                         std__mgr58__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane14_strm0_data        ;
  output                                        mgr58__std__lane14_strm0_data_valid  ;

  input                                         std__mgr58__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane14_strm1_data        ;
  output                                        mgr58__std__lane14_strm1_data_valid  ;

  input                                         std__mgr58__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane15_strm0_data        ;
  output                                        mgr58__std__lane15_strm0_data_valid  ;

  input                                         std__mgr58__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane15_strm1_data        ;
  output                                        mgr58__std__lane15_strm1_data_valid  ;

  input                                         std__mgr58__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane16_strm0_data        ;
  output                                        mgr58__std__lane16_strm0_data_valid  ;

  input                                         std__mgr58__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane16_strm1_data        ;
  output                                        mgr58__std__lane16_strm1_data_valid  ;

  input                                         std__mgr58__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane17_strm0_data        ;
  output                                        mgr58__std__lane17_strm0_data_valid  ;

  input                                         std__mgr58__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane17_strm1_data        ;
  output                                        mgr58__std__lane17_strm1_data_valid  ;

  input                                         std__mgr58__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane18_strm0_data        ;
  output                                        mgr58__std__lane18_strm0_data_valid  ;

  input                                         std__mgr58__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane18_strm1_data        ;
  output                                        mgr58__std__lane18_strm1_data_valid  ;

  input                                         std__mgr58__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane19_strm0_data        ;
  output                                        mgr58__std__lane19_strm0_data_valid  ;

  input                                         std__mgr58__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane19_strm1_data        ;
  output                                        mgr58__std__lane19_strm1_data_valid  ;

  input                                         std__mgr58__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane20_strm0_data        ;
  output                                        mgr58__std__lane20_strm0_data_valid  ;

  input                                         std__mgr58__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane20_strm1_data        ;
  output                                        mgr58__std__lane20_strm1_data_valid  ;

  input                                         std__mgr58__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane21_strm0_data        ;
  output                                        mgr58__std__lane21_strm0_data_valid  ;

  input                                         std__mgr58__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane21_strm1_data        ;
  output                                        mgr58__std__lane21_strm1_data_valid  ;

  input                                         std__mgr58__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane22_strm0_data        ;
  output                                        mgr58__std__lane22_strm0_data_valid  ;

  input                                         std__mgr58__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane22_strm1_data        ;
  output                                        mgr58__std__lane22_strm1_data_valid  ;

  input                                         std__mgr58__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane23_strm0_data        ;
  output                                        mgr58__std__lane23_strm0_data_valid  ;

  input                                         std__mgr58__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane23_strm1_data        ;
  output                                        mgr58__std__lane23_strm1_data_valid  ;

  input                                         std__mgr58__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane24_strm0_data        ;
  output                                        mgr58__std__lane24_strm0_data_valid  ;

  input                                         std__mgr58__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane24_strm1_data        ;
  output                                        mgr58__std__lane24_strm1_data_valid  ;

  input                                         std__mgr58__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane25_strm0_data        ;
  output                                        mgr58__std__lane25_strm0_data_valid  ;

  input                                         std__mgr58__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane25_strm1_data        ;
  output                                        mgr58__std__lane25_strm1_data_valid  ;

  input                                         std__mgr58__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane26_strm0_data        ;
  output                                        mgr58__std__lane26_strm0_data_valid  ;

  input                                         std__mgr58__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane26_strm1_data        ;
  output                                        mgr58__std__lane26_strm1_data_valid  ;

  input                                         std__mgr58__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane27_strm0_data        ;
  output                                        mgr58__std__lane27_strm0_data_valid  ;

  input                                         std__mgr58__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane27_strm1_data        ;
  output                                        mgr58__std__lane27_strm1_data_valid  ;

  input                                         std__mgr58__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane28_strm0_data        ;
  output                                        mgr58__std__lane28_strm0_data_valid  ;

  input                                         std__mgr58__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane28_strm1_data        ;
  output                                        mgr58__std__lane28_strm1_data_valid  ;

  input                                         std__mgr58__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane29_strm0_data        ;
  output                                        mgr58__std__lane29_strm0_data_valid  ;

  input                                         std__mgr58__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane29_strm1_data        ;
  output                                        mgr58__std__lane29_strm1_data_valid  ;

  input                                         std__mgr58__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane30_strm0_data        ;
  output                                        mgr58__std__lane30_strm0_data_valid  ;

  input                                         std__mgr58__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane30_strm1_data        ;
  output                                        mgr58__std__lane30_strm1_data_valid  ;

  input                                         std__mgr58__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane31_strm0_data        ;
  output                                        mgr58__std__lane31_strm0_data_valid  ;

  input                                         std__mgr58__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane31_strm1_data        ;
  output                                        mgr58__std__lane31_strm1_data_valid  ;

  input                                         std__mgr59__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane0_strm0_data        ;
  output                                        mgr59__std__lane0_strm0_data_valid  ;

  input                                         std__mgr59__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane0_strm1_data        ;
  output                                        mgr59__std__lane0_strm1_data_valid  ;

  input                                         std__mgr59__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane1_strm0_data        ;
  output                                        mgr59__std__lane1_strm0_data_valid  ;

  input                                         std__mgr59__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane1_strm1_data        ;
  output                                        mgr59__std__lane1_strm1_data_valid  ;

  input                                         std__mgr59__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane2_strm0_data        ;
  output                                        mgr59__std__lane2_strm0_data_valid  ;

  input                                         std__mgr59__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane2_strm1_data        ;
  output                                        mgr59__std__lane2_strm1_data_valid  ;

  input                                         std__mgr59__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane3_strm0_data        ;
  output                                        mgr59__std__lane3_strm0_data_valid  ;

  input                                         std__mgr59__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane3_strm1_data        ;
  output                                        mgr59__std__lane3_strm1_data_valid  ;

  input                                         std__mgr59__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane4_strm0_data        ;
  output                                        mgr59__std__lane4_strm0_data_valid  ;

  input                                         std__mgr59__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane4_strm1_data        ;
  output                                        mgr59__std__lane4_strm1_data_valid  ;

  input                                         std__mgr59__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane5_strm0_data        ;
  output                                        mgr59__std__lane5_strm0_data_valid  ;

  input                                         std__mgr59__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane5_strm1_data        ;
  output                                        mgr59__std__lane5_strm1_data_valid  ;

  input                                         std__mgr59__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane6_strm0_data        ;
  output                                        mgr59__std__lane6_strm0_data_valid  ;

  input                                         std__mgr59__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane6_strm1_data        ;
  output                                        mgr59__std__lane6_strm1_data_valid  ;

  input                                         std__mgr59__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane7_strm0_data        ;
  output                                        mgr59__std__lane7_strm0_data_valid  ;

  input                                         std__mgr59__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane7_strm1_data        ;
  output                                        mgr59__std__lane7_strm1_data_valid  ;

  input                                         std__mgr59__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane8_strm0_data        ;
  output                                        mgr59__std__lane8_strm0_data_valid  ;

  input                                         std__mgr59__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane8_strm1_data        ;
  output                                        mgr59__std__lane8_strm1_data_valid  ;

  input                                         std__mgr59__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane9_strm0_data        ;
  output                                        mgr59__std__lane9_strm0_data_valid  ;

  input                                         std__mgr59__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane9_strm1_data        ;
  output                                        mgr59__std__lane9_strm1_data_valid  ;

  input                                         std__mgr59__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane10_strm0_data        ;
  output                                        mgr59__std__lane10_strm0_data_valid  ;

  input                                         std__mgr59__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane10_strm1_data        ;
  output                                        mgr59__std__lane10_strm1_data_valid  ;

  input                                         std__mgr59__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane11_strm0_data        ;
  output                                        mgr59__std__lane11_strm0_data_valid  ;

  input                                         std__mgr59__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane11_strm1_data        ;
  output                                        mgr59__std__lane11_strm1_data_valid  ;

  input                                         std__mgr59__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane12_strm0_data        ;
  output                                        mgr59__std__lane12_strm0_data_valid  ;

  input                                         std__mgr59__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane12_strm1_data        ;
  output                                        mgr59__std__lane12_strm1_data_valid  ;

  input                                         std__mgr59__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane13_strm0_data        ;
  output                                        mgr59__std__lane13_strm0_data_valid  ;

  input                                         std__mgr59__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane13_strm1_data        ;
  output                                        mgr59__std__lane13_strm1_data_valid  ;

  input                                         std__mgr59__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane14_strm0_data        ;
  output                                        mgr59__std__lane14_strm0_data_valid  ;

  input                                         std__mgr59__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane14_strm1_data        ;
  output                                        mgr59__std__lane14_strm1_data_valid  ;

  input                                         std__mgr59__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane15_strm0_data        ;
  output                                        mgr59__std__lane15_strm0_data_valid  ;

  input                                         std__mgr59__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane15_strm1_data        ;
  output                                        mgr59__std__lane15_strm1_data_valid  ;

  input                                         std__mgr59__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane16_strm0_data        ;
  output                                        mgr59__std__lane16_strm0_data_valid  ;

  input                                         std__mgr59__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane16_strm1_data        ;
  output                                        mgr59__std__lane16_strm1_data_valid  ;

  input                                         std__mgr59__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane17_strm0_data        ;
  output                                        mgr59__std__lane17_strm0_data_valid  ;

  input                                         std__mgr59__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane17_strm1_data        ;
  output                                        mgr59__std__lane17_strm1_data_valid  ;

  input                                         std__mgr59__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane18_strm0_data        ;
  output                                        mgr59__std__lane18_strm0_data_valid  ;

  input                                         std__mgr59__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane18_strm1_data        ;
  output                                        mgr59__std__lane18_strm1_data_valid  ;

  input                                         std__mgr59__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane19_strm0_data        ;
  output                                        mgr59__std__lane19_strm0_data_valid  ;

  input                                         std__mgr59__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane19_strm1_data        ;
  output                                        mgr59__std__lane19_strm1_data_valid  ;

  input                                         std__mgr59__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane20_strm0_data        ;
  output                                        mgr59__std__lane20_strm0_data_valid  ;

  input                                         std__mgr59__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane20_strm1_data        ;
  output                                        mgr59__std__lane20_strm1_data_valid  ;

  input                                         std__mgr59__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane21_strm0_data        ;
  output                                        mgr59__std__lane21_strm0_data_valid  ;

  input                                         std__mgr59__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane21_strm1_data        ;
  output                                        mgr59__std__lane21_strm1_data_valid  ;

  input                                         std__mgr59__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane22_strm0_data        ;
  output                                        mgr59__std__lane22_strm0_data_valid  ;

  input                                         std__mgr59__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane22_strm1_data        ;
  output                                        mgr59__std__lane22_strm1_data_valid  ;

  input                                         std__mgr59__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane23_strm0_data        ;
  output                                        mgr59__std__lane23_strm0_data_valid  ;

  input                                         std__mgr59__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane23_strm1_data        ;
  output                                        mgr59__std__lane23_strm1_data_valid  ;

  input                                         std__mgr59__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane24_strm0_data        ;
  output                                        mgr59__std__lane24_strm0_data_valid  ;

  input                                         std__mgr59__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane24_strm1_data        ;
  output                                        mgr59__std__lane24_strm1_data_valid  ;

  input                                         std__mgr59__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane25_strm0_data        ;
  output                                        mgr59__std__lane25_strm0_data_valid  ;

  input                                         std__mgr59__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane25_strm1_data        ;
  output                                        mgr59__std__lane25_strm1_data_valid  ;

  input                                         std__mgr59__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane26_strm0_data        ;
  output                                        mgr59__std__lane26_strm0_data_valid  ;

  input                                         std__mgr59__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane26_strm1_data        ;
  output                                        mgr59__std__lane26_strm1_data_valid  ;

  input                                         std__mgr59__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane27_strm0_data        ;
  output                                        mgr59__std__lane27_strm0_data_valid  ;

  input                                         std__mgr59__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane27_strm1_data        ;
  output                                        mgr59__std__lane27_strm1_data_valid  ;

  input                                         std__mgr59__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane28_strm0_data        ;
  output                                        mgr59__std__lane28_strm0_data_valid  ;

  input                                         std__mgr59__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane28_strm1_data        ;
  output                                        mgr59__std__lane28_strm1_data_valid  ;

  input                                         std__mgr59__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane29_strm0_data        ;
  output                                        mgr59__std__lane29_strm0_data_valid  ;

  input                                         std__mgr59__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane29_strm1_data        ;
  output                                        mgr59__std__lane29_strm1_data_valid  ;

  input                                         std__mgr59__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane30_strm0_data        ;
  output                                        mgr59__std__lane30_strm0_data_valid  ;

  input                                         std__mgr59__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane30_strm1_data        ;
  output                                        mgr59__std__lane30_strm1_data_valid  ;

  input                                         std__mgr59__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane31_strm0_data        ;
  output                                        mgr59__std__lane31_strm0_data_valid  ;

  input                                         std__mgr59__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane31_strm1_data        ;
  output                                        mgr59__std__lane31_strm1_data_valid  ;

  input                                         std__mgr60__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane0_strm0_data        ;
  output                                        mgr60__std__lane0_strm0_data_valid  ;

  input                                         std__mgr60__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane0_strm1_data        ;
  output                                        mgr60__std__lane0_strm1_data_valid  ;

  input                                         std__mgr60__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane1_strm0_data        ;
  output                                        mgr60__std__lane1_strm0_data_valid  ;

  input                                         std__mgr60__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane1_strm1_data        ;
  output                                        mgr60__std__lane1_strm1_data_valid  ;

  input                                         std__mgr60__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane2_strm0_data        ;
  output                                        mgr60__std__lane2_strm0_data_valid  ;

  input                                         std__mgr60__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane2_strm1_data        ;
  output                                        mgr60__std__lane2_strm1_data_valid  ;

  input                                         std__mgr60__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane3_strm0_data        ;
  output                                        mgr60__std__lane3_strm0_data_valid  ;

  input                                         std__mgr60__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane3_strm1_data        ;
  output                                        mgr60__std__lane3_strm1_data_valid  ;

  input                                         std__mgr60__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane4_strm0_data        ;
  output                                        mgr60__std__lane4_strm0_data_valid  ;

  input                                         std__mgr60__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane4_strm1_data        ;
  output                                        mgr60__std__lane4_strm1_data_valid  ;

  input                                         std__mgr60__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane5_strm0_data        ;
  output                                        mgr60__std__lane5_strm0_data_valid  ;

  input                                         std__mgr60__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane5_strm1_data        ;
  output                                        mgr60__std__lane5_strm1_data_valid  ;

  input                                         std__mgr60__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane6_strm0_data        ;
  output                                        mgr60__std__lane6_strm0_data_valid  ;

  input                                         std__mgr60__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane6_strm1_data        ;
  output                                        mgr60__std__lane6_strm1_data_valid  ;

  input                                         std__mgr60__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane7_strm0_data        ;
  output                                        mgr60__std__lane7_strm0_data_valid  ;

  input                                         std__mgr60__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane7_strm1_data        ;
  output                                        mgr60__std__lane7_strm1_data_valid  ;

  input                                         std__mgr60__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane8_strm0_data        ;
  output                                        mgr60__std__lane8_strm0_data_valid  ;

  input                                         std__mgr60__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane8_strm1_data        ;
  output                                        mgr60__std__lane8_strm1_data_valid  ;

  input                                         std__mgr60__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane9_strm0_data        ;
  output                                        mgr60__std__lane9_strm0_data_valid  ;

  input                                         std__mgr60__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane9_strm1_data        ;
  output                                        mgr60__std__lane9_strm1_data_valid  ;

  input                                         std__mgr60__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane10_strm0_data        ;
  output                                        mgr60__std__lane10_strm0_data_valid  ;

  input                                         std__mgr60__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane10_strm1_data        ;
  output                                        mgr60__std__lane10_strm1_data_valid  ;

  input                                         std__mgr60__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane11_strm0_data        ;
  output                                        mgr60__std__lane11_strm0_data_valid  ;

  input                                         std__mgr60__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane11_strm1_data        ;
  output                                        mgr60__std__lane11_strm1_data_valid  ;

  input                                         std__mgr60__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane12_strm0_data        ;
  output                                        mgr60__std__lane12_strm0_data_valid  ;

  input                                         std__mgr60__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane12_strm1_data        ;
  output                                        mgr60__std__lane12_strm1_data_valid  ;

  input                                         std__mgr60__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane13_strm0_data        ;
  output                                        mgr60__std__lane13_strm0_data_valid  ;

  input                                         std__mgr60__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane13_strm1_data        ;
  output                                        mgr60__std__lane13_strm1_data_valid  ;

  input                                         std__mgr60__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane14_strm0_data        ;
  output                                        mgr60__std__lane14_strm0_data_valid  ;

  input                                         std__mgr60__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane14_strm1_data        ;
  output                                        mgr60__std__lane14_strm1_data_valid  ;

  input                                         std__mgr60__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane15_strm0_data        ;
  output                                        mgr60__std__lane15_strm0_data_valid  ;

  input                                         std__mgr60__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane15_strm1_data        ;
  output                                        mgr60__std__lane15_strm1_data_valid  ;

  input                                         std__mgr60__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane16_strm0_data        ;
  output                                        mgr60__std__lane16_strm0_data_valid  ;

  input                                         std__mgr60__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane16_strm1_data        ;
  output                                        mgr60__std__lane16_strm1_data_valid  ;

  input                                         std__mgr60__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane17_strm0_data        ;
  output                                        mgr60__std__lane17_strm0_data_valid  ;

  input                                         std__mgr60__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane17_strm1_data        ;
  output                                        mgr60__std__lane17_strm1_data_valid  ;

  input                                         std__mgr60__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane18_strm0_data        ;
  output                                        mgr60__std__lane18_strm0_data_valid  ;

  input                                         std__mgr60__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane18_strm1_data        ;
  output                                        mgr60__std__lane18_strm1_data_valid  ;

  input                                         std__mgr60__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane19_strm0_data        ;
  output                                        mgr60__std__lane19_strm0_data_valid  ;

  input                                         std__mgr60__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane19_strm1_data        ;
  output                                        mgr60__std__lane19_strm1_data_valid  ;

  input                                         std__mgr60__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane20_strm0_data        ;
  output                                        mgr60__std__lane20_strm0_data_valid  ;

  input                                         std__mgr60__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane20_strm1_data        ;
  output                                        mgr60__std__lane20_strm1_data_valid  ;

  input                                         std__mgr60__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane21_strm0_data        ;
  output                                        mgr60__std__lane21_strm0_data_valid  ;

  input                                         std__mgr60__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane21_strm1_data        ;
  output                                        mgr60__std__lane21_strm1_data_valid  ;

  input                                         std__mgr60__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane22_strm0_data        ;
  output                                        mgr60__std__lane22_strm0_data_valid  ;

  input                                         std__mgr60__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane22_strm1_data        ;
  output                                        mgr60__std__lane22_strm1_data_valid  ;

  input                                         std__mgr60__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane23_strm0_data        ;
  output                                        mgr60__std__lane23_strm0_data_valid  ;

  input                                         std__mgr60__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane23_strm1_data        ;
  output                                        mgr60__std__lane23_strm1_data_valid  ;

  input                                         std__mgr60__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane24_strm0_data        ;
  output                                        mgr60__std__lane24_strm0_data_valid  ;

  input                                         std__mgr60__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane24_strm1_data        ;
  output                                        mgr60__std__lane24_strm1_data_valid  ;

  input                                         std__mgr60__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane25_strm0_data        ;
  output                                        mgr60__std__lane25_strm0_data_valid  ;

  input                                         std__mgr60__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane25_strm1_data        ;
  output                                        mgr60__std__lane25_strm1_data_valid  ;

  input                                         std__mgr60__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane26_strm0_data        ;
  output                                        mgr60__std__lane26_strm0_data_valid  ;

  input                                         std__mgr60__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane26_strm1_data        ;
  output                                        mgr60__std__lane26_strm1_data_valid  ;

  input                                         std__mgr60__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane27_strm0_data        ;
  output                                        mgr60__std__lane27_strm0_data_valid  ;

  input                                         std__mgr60__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane27_strm1_data        ;
  output                                        mgr60__std__lane27_strm1_data_valid  ;

  input                                         std__mgr60__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane28_strm0_data        ;
  output                                        mgr60__std__lane28_strm0_data_valid  ;

  input                                         std__mgr60__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane28_strm1_data        ;
  output                                        mgr60__std__lane28_strm1_data_valid  ;

  input                                         std__mgr60__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane29_strm0_data        ;
  output                                        mgr60__std__lane29_strm0_data_valid  ;

  input                                         std__mgr60__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane29_strm1_data        ;
  output                                        mgr60__std__lane29_strm1_data_valid  ;

  input                                         std__mgr60__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane30_strm0_data        ;
  output                                        mgr60__std__lane30_strm0_data_valid  ;

  input                                         std__mgr60__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane30_strm1_data        ;
  output                                        mgr60__std__lane30_strm1_data_valid  ;

  input                                         std__mgr60__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane31_strm0_data        ;
  output                                        mgr60__std__lane31_strm0_data_valid  ;

  input                                         std__mgr60__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane31_strm1_data        ;
  output                                        mgr60__std__lane31_strm1_data_valid  ;

  input                                         std__mgr61__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane0_strm0_data        ;
  output                                        mgr61__std__lane0_strm0_data_valid  ;

  input                                         std__mgr61__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane0_strm1_data        ;
  output                                        mgr61__std__lane0_strm1_data_valid  ;

  input                                         std__mgr61__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane1_strm0_data        ;
  output                                        mgr61__std__lane1_strm0_data_valid  ;

  input                                         std__mgr61__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane1_strm1_data        ;
  output                                        mgr61__std__lane1_strm1_data_valid  ;

  input                                         std__mgr61__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane2_strm0_data        ;
  output                                        mgr61__std__lane2_strm0_data_valid  ;

  input                                         std__mgr61__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane2_strm1_data        ;
  output                                        mgr61__std__lane2_strm1_data_valid  ;

  input                                         std__mgr61__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane3_strm0_data        ;
  output                                        mgr61__std__lane3_strm0_data_valid  ;

  input                                         std__mgr61__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane3_strm1_data        ;
  output                                        mgr61__std__lane3_strm1_data_valid  ;

  input                                         std__mgr61__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane4_strm0_data        ;
  output                                        mgr61__std__lane4_strm0_data_valid  ;

  input                                         std__mgr61__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane4_strm1_data        ;
  output                                        mgr61__std__lane4_strm1_data_valid  ;

  input                                         std__mgr61__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane5_strm0_data        ;
  output                                        mgr61__std__lane5_strm0_data_valid  ;

  input                                         std__mgr61__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane5_strm1_data        ;
  output                                        mgr61__std__lane5_strm1_data_valid  ;

  input                                         std__mgr61__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane6_strm0_data        ;
  output                                        mgr61__std__lane6_strm0_data_valid  ;

  input                                         std__mgr61__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane6_strm1_data        ;
  output                                        mgr61__std__lane6_strm1_data_valid  ;

  input                                         std__mgr61__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane7_strm0_data        ;
  output                                        mgr61__std__lane7_strm0_data_valid  ;

  input                                         std__mgr61__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane7_strm1_data        ;
  output                                        mgr61__std__lane7_strm1_data_valid  ;

  input                                         std__mgr61__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane8_strm0_data        ;
  output                                        mgr61__std__lane8_strm0_data_valid  ;

  input                                         std__mgr61__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane8_strm1_data        ;
  output                                        mgr61__std__lane8_strm1_data_valid  ;

  input                                         std__mgr61__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane9_strm0_data        ;
  output                                        mgr61__std__lane9_strm0_data_valid  ;

  input                                         std__mgr61__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane9_strm1_data        ;
  output                                        mgr61__std__lane9_strm1_data_valid  ;

  input                                         std__mgr61__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane10_strm0_data        ;
  output                                        mgr61__std__lane10_strm0_data_valid  ;

  input                                         std__mgr61__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane10_strm1_data        ;
  output                                        mgr61__std__lane10_strm1_data_valid  ;

  input                                         std__mgr61__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane11_strm0_data        ;
  output                                        mgr61__std__lane11_strm0_data_valid  ;

  input                                         std__mgr61__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane11_strm1_data        ;
  output                                        mgr61__std__lane11_strm1_data_valid  ;

  input                                         std__mgr61__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane12_strm0_data        ;
  output                                        mgr61__std__lane12_strm0_data_valid  ;

  input                                         std__mgr61__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane12_strm1_data        ;
  output                                        mgr61__std__lane12_strm1_data_valid  ;

  input                                         std__mgr61__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane13_strm0_data        ;
  output                                        mgr61__std__lane13_strm0_data_valid  ;

  input                                         std__mgr61__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane13_strm1_data        ;
  output                                        mgr61__std__lane13_strm1_data_valid  ;

  input                                         std__mgr61__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane14_strm0_data        ;
  output                                        mgr61__std__lane14_strm0_data_valid  ;

  input                                         std__mgr61__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane14_strm1_data        ;
  output                                        mgr61__std__lane14_strm1_data_valid  ;

  input                                         std__mgr61__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane15_strm0_data        ;
  output                                        mgr61__std__lane15_strm0_data_valid  ;

  input                                         std__mgr61__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane15_strm1_data        ;
  output                                        mgr61__std__lane15_strm1_data_valid  ;

  input                                         std__mgr61__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane16_strm0_data        ;
  output                                        mgr61__std__lane16_strm0_data_valid  ;

  input                                         std__mgr61__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane16_strm1_data        ;
  output                                        mgr61__std__lane16_strm1_data_valid  ;

  input                                         std__mgr61__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane17_strm0_data        ;
  output                                        mgr61__std__lane17_strm0_data_valid  ;

  input                                         std__mgr61__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane17_strm1_data        ;
  output                                        mgr61__std__lane17_strm1_data_valid  ;

  input                                         std__mgr61__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane18_strm0_data        ;
  output                                        mgr61__std__lane18_strm0_data_valid  ;

  input                                         std__mgr61__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane18_strm1_data        ;
  output                                        mgr61__std__lane18_strm1_data_valid  ;

  input                                         std__mgr61__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane19_strm0_data        ;
  output                                        mgr61__std__lane19_strm0_data_valid  ;

  input                                         std__mgr61__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane19_strm1_data        ;
  output                                        mgr61__std__lane19_strm1_data_valid  ;

  input                                         std__mgr61__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane20_strm0_data        ;
  output                                        mgr61__std__lane20_strm0_data_valid  ;

  input                                         std__mgr61__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane20_strm1_data        ;
  output                                        mgr61__std__lane20_strm1_data_valid  ;

  input                                         std__mgr61__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane21_strm0_data        ;
  output                                        mgr61__std__lane21_strm0_data_valid  ;

  input                                         std__mgr61__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane21_strm1_data        ;
  output                                        mgr61__std__lane21_strm1_data_valid  ;

  input                                         std__mgr61__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane22_strm0_data        ;
  output                                        mgr61__std__lane22_strm0_data_valid  ;

  input                                         std__mgr61__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane22_strm1_data        ;
  output                                        mgr61__std__lane22_strm1_data_valid  ;

  input                                         std__mgr61__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane23_strm0_data        ;
  output                                        mgr61__std__lane23_strm0_data_valid  ;

  input                                         std__mgr61__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane23_strm1_data        ;
  output                                        mgr61__std__lane23_strm1_data_valid  ;

  input                                         std__mgr61__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane24_strm0_data        ;
  output                                        mgr61__std__lane24_strm0_data_valid  ;

  input                                         std__mgr61__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane24_strm1_data        ;
  output                                        mgr61__std__lane24_strm1_data_valid  ;

  input                                         std__mgr61__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane25_strm0_data        ;
  output                                        mgr61__std__lane25_strm0_data_valid  ;

  input                                         std__mgr61__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane25_strm1_data        ;
  output                                        mgr61__std__lane25_strm1_data_valid  ;

  input                                         std__mgr61__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane26_strm0_data        ;
  output                                        mgr61__std__lane26_strm0_data_valid  ;

  input                                         std__mgr61__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane26_strm1_data        ;
  output                                        mgr61__std__lane26_strm1_data_valid  ;

  input                                         std__mgr61__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane27_strm0_data        ;
  output                                        mgr61__std__lane27_strm0_data_valid  ;

  input                                         std__mgr61__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane27_strm1_data        ;
  output                                        mgr61__std__lane27_strm1_data_valid  ;

  input                                         std__mgr61__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane28_strm0_data        ;
  output                                        mgr61__std__lane28_strm0_data_valid  ;

  input                                         std__mgr61__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane28_strm1_data        ;
  output                                        mgr61__std__lane28_strm1_data_valid  ;

  input                                         std__mgr61__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane29_strm0_data        ;
  output                                        mgr61__std__lane29_strm0_data_valid  ;

  input                                         std__mgr61__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane29_strm1_data        ;
  output                                        mgr61__std__lane29_strm1_data_valid  ;

  input                                         std__mgr61__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane30_strm0_data        ;
  output                                        mgr61__std__lane30_strm0_data_valid  ;

  input                                         std__mgr61__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane30_strm1_data        ;
  output                                        mgr61__std__lane30_strm1_data_valid  ;

  input                                         std__mgr61__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane31_strm0_data        ;
  output                                        mgr61__std__lane31_strm0_data_valid  ;

  input                                         std__mgr61__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane31_strm1_data        ;
  output                                        mgr61__std__lane31_strm1_data_valid  ;

  input                                         std__mgr62__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane0_strm0_data        ;
  output                                        mgr62__std__lane0_strm0_data_valid  ;

  input                                         std__mgr62__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane0_strm1_data        ;
  output                                        mgr62__std__lane0_strm1_data_valid  ;

  input                                         std__mgr62__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane1_strm0_data        ;
  output                                        mgr62__std__lane1_strm0_data_valid  ;

  input                                         std__mgr62__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane1_strm1_data        ;
  output                                        mgr62__std__lane1_strm1_data_valid  ;

  input                                         std__mgr62__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane2_strm0_data        ;
  output                                        mgr62__std__lane2_strm0_data_valid  ;

  input                                         std__mgr62__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane2_strm1_data        ;
  output                                        mgr62__std__lane2_strm1_data_valid  ;

  input                                         std__mgr62__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane3_strm0_data        ;
  output                                        mgr62__std__lane3_strm0_data_valid  ;

  input                                         std__mgr62__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane3_strm1_data        ;
  output                                        mgr62__std__lane3_strm1_data_valid  ;

  input                                         std__mgr62__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane4_strm0_data        ;
  output                                        mgr62__std__lane4_strm0_data_valid  ;

  input                                         std__mgr62__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane4_strm1_data        ;
  output                                        mgr62__std__lane4_strm1_data_valid  ;

  input                                         std__mgr62__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane5_strm0_data        ;
  output                                        mgr62__std__lane5_strm0_data_valid  ;

  input                                         std__mgr62__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane5_strm1_data        ;
  output                                        mgr62__std__lane5_strm1_data_valid  ;

  input                                         std__mgr62__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane6_strm0_data        ;
  output                                        mgr62__std__lane6_strm0_data_valid  ;

  input                                         std__mgr62__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane6_strm1_data        ;
  output                                        mgr62__std__lane6_strm1_data_valid  ;

  input                                         std__mgr62__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane7_strm0_data        ;
  output                                        mgr62__std__lane7_strm0_data_valid  ;

  input                                         std__mgr62__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane7_strm1_data        ;
  output                                        mgr62__std__lane7_strm1_data_valid  ;

  input                                         std__mgr62__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane8_strm0_data        ;
  output                                        mgr62__std__lane8_strm0_data_valid  ;

  input                                         std__mgr62__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane8_strm1_data        ;
  output                                        mgr62__std__lane8_strm1_data_valid  ;

  input                                         std__mgr62__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane9_strm0_data        ;
  output                                        mgr62__std__lane9_strm0_data_valid  ;

  input                                         std__mgr62__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane9_strm1_data        ;
  output                                        mgr62__std__lane9_strm1_data_valid  ;

  input                                         std__mgr62__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane10_strm0_data        ;
  output                                        mgr62__std__lane10_strm0_data_valid  ;

  input                                         std__mgr62__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane10_strm1_data        ;
  output                                        mgr62__std__lane10_strm1_data_valid  ;

  input                                         std__mgr62__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane11_strm0_data        ;
  output                                        mgr62__std__lane11_strm0_data_valid  ;

  input                                         std__mgr62__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane11_strm1_data        ;
  output                                        mgr62__std__lane11_strm1_data_valid  ;

  input                                         std__mgr62__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane12_strm0_data        ;
  output                                        mgr62__std__lane12_strm0_data_valid  ;

  input                                         std__mgr62__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane12_strm1_data        ;
  output                                        mgr62__std__lane12_strm1_data_valid  ;

  input                                         std__mgr62__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane13_strm0_data        ;
  output                                        mgr62__std__lane13_strm0_data_valid  ;

  input                                         std__mgr62__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane13_strm1_data        ;
  output                                        mgr62__std__lane13_strm1_data_valid  ;

  input                                         std__mgr62__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane14_strm0_data        ;
  output                                        mgr62__std__lane14_strm0_data_valid  ;

  input                                         std__mgr62__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane14_strm1_data        ;
  output                                        mgr62__std__lane14_strm1_data_valid  ;

  input                                         std__mgr62__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane15_strm0_data        ;
  output                                        mgr62__std__lane15_strm0_data_valid  ;

  input                                         std__mgr62__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane15_strm1_data        ;
  output                                        mgr62__std__lane15_strm1_data_valid  ;

  input                                         std__mgr62__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane16_strm0_data        ;
  output                                        mgr62__std__lane16_strm0_data_valid  ;

  input                                         std__mgr62__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane16_strm1_data        ;
  output                                        mgr62__std__lane16_strm1_data_valid  ;

  input                                         std__mgr62__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane17_strm0_data        ;
  output                                        mgr62__std__lane17_strm0_data_valid  ;

  input                                         std__mgr62__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane17_strm1_data        ;
  output                                        mgr62__std__lane17_strm1_data_valid  ;

  input                                         std__mgr62__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane18_strm0_data        ;
  output                                        mgr62__std__lane18_strm0_data_valid  ;

  input                                         std__mgr62__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane18_strm1_data        ;
  output                                        mgr62__std__lane18_strm1_data_valid  ;

  input                                         std__mgr62__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane19_strm0_data        ;
  output                                        mgr62__std__lane19_strm0_data_valid  ;

  input                                         std__mgr62__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane19_strm1_data        ;
  output                                        mgr62__std__lane19_strm1_data_valid  ;

  input                                         std__mgr62__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane20_strm0_data        ;
  output                                        mgr62__std__lane20_strm0_data_valid  ;

  input                                         std__mgr62__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane20_strm1_data        ;
  output                                        mgr62__std__lane20_strm1_data_valid  ;

  input                                         std__mgr62__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane21_strm0_data        ;
  output                                        mgr62__std__lane21_strm0_data_valid  ;

  input                                         std__mgr62__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane21_strm1_data        ;
  output                                        mgr62__std__lane21_strm1_data_valid  ;

  input                                         std__mgr62__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane22_strm0_data        ;
  output                                        mgr62__std__lane22_strm0_data_valid  ;

  input                                         std__mgr62__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane22_strm1_data        ;
  output                                        mgr62__std__lane22_strm1_data_valid  ;

  input                                         std__mgr62__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane23_strm0_data        ;
  output                                        mgr62__std__lane23_strm0_data_valid  ;

  input                                         std__mgr62__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane23_strm1_data        ;
  output                                        mgr62__std__lane23_strm1_data_valid  ;

  input                                         std__mgr62__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane24_strm0_data        ;
  output                                        mgr62__std__lane24_strm0_data_valid  ;

  input                                         std__mgr62__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane24_strm1_data        ;
  output                                        mgr62__std__lane24_strm1_data_valid  ;

  input                                         std__mgr62__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane25_strm0_data        ;
  output                                        mgr62__std__lane25_strm0_data_valid  ;

  input                                         std__mgr62__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane25_strm1_data        ;
  output                                        mgr62__std__lane25_strm1_data_valid  ;

  input                                         std__mgr62__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane26_strm0_data        ;
  output                                        mgr62__std__lane26_strm0_data_valid  ;

  input                                         std__mgr62__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane26_strm1_data        ;
  output                                        mgr62__std__lane26_strm1_data_valid  ;

  input                                         std__mgr62__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane27_strm0_data        ;
  output                                        mgr62__std__lane27_strm0_data_valid  ;

  input                                         std__mgr62__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane27_strm1_data        ;
  output                                        mgr62__std__lane27_strm1_data_valid  ;

  input                                         std__mgr62__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane28_strm0_data        ;
  output                                        mgr62__std__lane28_strm0_data_valid  ;

  input                                         std__mgr62__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane28_strm1_data        ;
  output                                        mgr62__std__lane28_strm1_data_valid  ;

  input                                         std__mgr62__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane29_strm0_data        ;
  output                                        mgr62__std__lane29_strm0_data_valid  ;

  input                                         std__mgr62__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane29_strm1_data        ;
  output                                        mgr62__std__lane29_strm1_data_valid  ;

  input                                         std__mgr62__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane30_strm0_data        ;
  output                                        mgr62__std__lane30_strm0_data_valid  ;

  input                                         std__mgr62__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane30_strm1_data        ;
  output                                        mgr62__std__lane30_strm1_data_valid  ;

  input                                         std__mgr62__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane31_strm0_data        ;
  output                                        mgr62__std__lane31_strm0_data_valid  ;

  input                                         std__mgr62__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane31_strm1_data        ;
  output                                        mgr62__std__lane31_strm1_data_valid  ;

  input                                         std__mgr63__lane0_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane0_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane0_strm0_data        ;
  output                                        mgr63__std__lane0_strm0_data_valid  ;

  input                                         std__mgr63__lane0_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane0_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane0_strm1_data        ;
  output                                        mgr63__std__lane0_strm1_data_valid  ;

  input                                         std__mgr63__lane1_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane1_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane1_strm0_data        ;
  output                                        mgr63__std__lane1_strm0_data_valid  ;

  input                                         std__mgr63__lane1_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane1_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane1_strm1_data        ;
  output                                        mgr63__std__lane1_strm1_data_valid  ;

  input                                         std__mgr63__lane2_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane2_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane2_strm0_data        ;
  output                                        mgr63__std__lane2_strm0_data_valid  ;

  input                                         std__mgr63__lane2_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane2_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane2_strm1_data        ;
  output                                        mgr63__std__lane2_strm1_data_valid  ;

  input                                         std__mgr63__lane3_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane3_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane3_strm0_data        ;
  output                                        mgr63__std__lane3_strm0_data_valid  ;

  input                                         std__mgr63__lane3_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane3_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane3_strm1_data        ;
  output                                        mgr63__std__lane3_strm1_data_valid  ;

  input                                         std__mgr63__lane4_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane4_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane4_strm0_data        ;
  output                                        mgr63__std__lane4_strm0_data_valid  ;

  input                                         std__mgr63__lane4_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane4_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane4_strm1_data        ;
  output                                        mgr63__std__lane4_strm1_data_valid  ;

  input                                         std__mgr63__lane5_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane5_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane5_strm0_data        ;
  output                                        mgr63__std__lane5_strm0_data_valid  ;

  input                                         std__mgr63__lane5_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane5_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane5_strm1_data        ;
  output                                        mgr63__std__lane5_strm1_data_valid  ;

  input                                         std__mgr63__lane6_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane6_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane6_strm0_data        ;
  output                                        mgr63__std__lane6_strm0_data_valid  ;

  input                                         std__mgr63__lane6_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane6_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane6_strm1_data        ;
  output                                        mgr63__std__lane6_strm1_data_valid  ;

  input                                         std__mgr63__lane7_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane7_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane7_strm0_data        ;
  output                                        mgr63__std__lane7_strm0_data_valid  ;

  input                                         std__mgr63__lane7_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane7_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane7_strm1_data        ;
  output                                        mgr63__std__lane7_strm1_data_valid  ;

  input                                         std__mgr63__lane8_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane8_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane8_strm0_data        ;
  output                                        mgr63__std__lane8_strm0_data_valid  ;

  input                                         std__mgr63__lane8_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane8_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane8_strm1_data        ;
  output                                        mgr63__std__lane8_strm1_data_valid  ;

  input                                         std__mgr63__lane9_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane9_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane9_strm0_data        ;
  output                                        mgr63__std__lane9_strm0_data_valid  ;

  input                                         std__mgr63__lane9_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane9_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane9_strm1_data        ;
  output                                        mgr63__std__lane9_strm1_data_valid  ;

  input                                         std__mgr63__lane10_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane10_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane10_strm0_data        ;
  output                                        mgr63__std__lane10_strm0_data_valid  ;

  input                                         std__mgr63__lane10_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane10_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane10_strm1_data        ;
  output                                        mgr63__std__lane10_strm1_data_valid  ;

  input                                         std__mgr63__lane11_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane11_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane11_strm0_data        ;
  output                                        mgr63__std__lane11_strm0_data_valid  ;

  input                                         std__mgr63__lane11_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane11_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane11_strm1_data        ;
  output                                        mgr63__std__lane11_strm1_data_valid  ;

  input                                         std__mgr63__lane12_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane12_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane12_strm0_data        ;
  output                                        mgr63__std__lane12_strm0_data_valid  ;

  input                                         std__mgr63__lane12_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane12_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane12_strm1_data        ;
  output                                        mgr63__std__lane12_strm1_data_valid  ;

  input                                         std__mgr63__lane13_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane13_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane13_strm0_data        ;
  output                                        mgr63__std__lane13_strm0_data_valid  ;

  input                                         std__mgr63__lane13_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane13_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane13_strm1_data        ;
  output                                        mgr63__std__lane13_strm1_data_valid  ;

  input                                         std__mgr63__lane14_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane14_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane14_strm0_data        ;
  output                                        mgr63__std__lane14_strm0_data_valid  ;

  input                                         std__mgr63__lane14_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane14_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane14_strm1_data        ;
  output                                        mgr63__std__lane14_strm1_data_valid  ;

  input                                         std__mgr63__lane15_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane15_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane15_strm0_data        ;
  output                                        mgr63__std__lane15_strm0_data_valid  ;

  input                                         std__mgr63__lane15_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane15_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane15_strm1_data        ;
  output                                        mgr63__std__lane15_strm1_data_valid  ;

  input                                         std__mgr63__lane16_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane16_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane16_strm0_data        ;
  output                                        mgr63__std__lane16_strm0_data_valid  ;

  input                                         std__mgr63__lane16_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane16_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane16_strm1_data        ;
  output                                        mgr63__std__lane16_strm1_data_valid  ;

  input                                         std__mgr63__lane17_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane17_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane17_strm0_data        ;
  output                                        mgr63__std__lane17_strm0_data_valid  ;

  input                                         std__mgr63__lane17_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane17_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane17_strm1_data        ;
  output                                        mgr63__std__lane17_strm1_data_valid  ;

  input                                         std__mgr63__lane18_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane18_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane18_strm0_data        ;
  output                                        mgr63__std__lane18_strm0_data_valid  ;

  input                                         std__mgr63__lane18_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane18_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane18_strm1_data        ;
  output                                        mgr63__std__lane18_strm1_data_valid  ;

  input                                         std__mgr63__lane19_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane19_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane19_strm0_data        ;
  output                                        mgr63__std__lane19_strm0_data_valid  ;

  input                                         std__mgr63__lane19_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane19_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane19_strm1_data        ;
  output                                        mgr63__std__lane19_strm1_data_valid  ;

  input                                         std__mgr63__lane20_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane20_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane20_strm0_data        ;
  output                                        mgr63__std__lane20_strm0_data_valid  ;

  input                                         std__mgr63__lane20_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane20_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane20_strm1_data        ;
  output                                        mgr63__std__lane20_strm1_data_valid  ;

  input                                         std__mgr63__lane21_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane21_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane21_strm0_data        ;
  output                                        mgr63__std__lane21_strm0_data_valid  ;

  input                                         std__mgr63__lane21_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane21_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane21_strm1_data        ;
  output                                        mgr63__std__lane21_strm1_data_valid  ;

  input                                         std__mgr63__lane22_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane22_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane22_strm0_data        ;
  output                                        mgr63__std__lane22_strm0_data_valid  ;

  input                                         std__mgr63__lane22_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane22_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane22_strm1_data        ;
  output                                        mgr63__std__lane22_strm1_data_valid  ;

  input                                         std__mgr63__lane23_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane23_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane23_strm0_data        ;
  output                                        mgr63__std__lane23_strm0_data_valid  ;

  input                                         std__mgr63__lane23_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane23_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane23_strm1_data        ;
  output                                        mgr63__std__lane23_strm1_data_valid  ;

  input                                         std__mgr63__lane24_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane24_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane24_strm0_data        ;
  output                                        mgr63__std__lane24_strm0_data_valid  ;

  input                                         std__mgr63__lane24_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane24_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane24_strm1_data        ;
  output                                        mgr63__std__lane24_strm1_data_valid  ;

  input                                         std__mgr63__lane25_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane25_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane25_strm0_data        ;
  output                                        mgr63__std__lane25_strm0_data_valid  ;

  input                                         std__mgr63__lane25_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane25_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane25_strm1_data        ;
  output                                        mgr63__std__lane25_strm1_data_valid  ;

  input                                         std__mgr63__lane26_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane26_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane26_strm0_data        ;
  output                                        mgr63__std__lane26_strm0_data_valid  ;

  input                                         std__mgr63__lane26_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane26_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane26_strm1_data        ;
  output                                        mgr63__std__lane26_strm1_data_valid  ;

  input                                         std__mgr63__lane27_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane27_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane27_strm0_data        ;
  output                                        mgr63__std__lane27_strm0_data_valid  ;

  input                                         std__mgr63__lane27_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane27_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane27_strm1_data        ;
  output                                        mgr63__std__lane27_strm1_data_valid  ;

  input                                         std__mgr63__lane28_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane28_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane28_strm0_data        ;
  output                                        mgr63__std__lane28_strm0_data_valid  ;

  input                                         std__mgr63__lane28_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane28_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane28_strm1_data        ;
  output                                        mgr63__std__lane28_strm1_data_valid  ;

  input                                         std__mgr63__lane29_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane29_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane29_strm0_data        ;
  output                                        mgr63__std__lane29_strm0_data_valid  ;

  input                                         std__mgr63__lane29_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane29_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane29_strm1_data        ;
  output                                        mgr63__std__lane29_strm1_data_valid  ;

  input                                         std__mgr63__lane30_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane30_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane30_strm0_data        ;
  output                                        mgr63__std__lane30_strm0_data_valid  ;

  input                                         std__mgr63__lane30_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane30_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane30_strm1_data        ;
  output                                        mgr63__std__lane30_strm1_data_valid  ;

  input                                         std__mgr63__lane31_strm0_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane31_strm0_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane31_strm0_data        ;
  output                                        mgr63__std__lane31_strm0_data_valid  ;

  input                                         std__mgr63__lane31_strm1_ready       ;
  output  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane31_strm1_cntl        ;
  output  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane31_strm1_data        ;
  output                                        mgr63__std__lane31_strm1_data_valid  ;
