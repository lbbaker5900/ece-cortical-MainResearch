
  // General control and status                                                   
  output                                        mgr0__sys__allSynchronized     ;
  input                                         sys__mgr0__thisSynchronized    ;
  input                                         sys__mgr0__ready               ;
  input                                         sys__mgr0__complete            ;
  // General control and status                                                   
  output                                        mgr1__sys__allSynchronized     ;
  input                                         sys__mgr1__thisSynchronized    ;
  input                                         sys__mgr1__ready               ;
  input                                         sys__mgr1__complete            ;
  // General control and status                                                   
  output                                        mgr2__sys__allSynchronized     ;
  input                                         sys__mgr2__thisSynchronized    ;
  input                                         sys__mgr2__ready               ;
  input                                         sys__mgr2__complete            ;
  // General control and status                                                   
  output                                        mgr3__sys__allSynchronized     ;
  input                                         sys__mgr3__thisSynchronized    ;
  input                                         sys__mgr3__ready               ;
  input                                         sys__mgr3__complete            ;
  // General control and status                                                   
  output                                        mgr4__sys__allSynchronized     ;
  input                                         sys__mgr4__thisSynchronized    ;
  input                                         sys__mgr4__ready               ;
  input                                         sys__mgr4__complete            ;
  // General control and status                                                   
  output                                        mgr5__sys__allSynchronized     ;
  input                                         sys__mgr5__thisSynchronized    ;
  input                                         sys__mgr5__ready               ;
  input                                         sys__mgr5__complete            ;
  // General control and status                                                   
  output                                        mgr6__sys__allSynchronized     ;
  input                                         sys__mgr6__thisSynchronized    ;
  input                                         sys__mgr6__ready               ;
  input                                         sys__mgr6__complete            ;
  // General control and status                                                   
  output                                        mgr7__sys__allSynchronized     ;
  input                                         sys__mgr7__thisSynchronized    ;
  input                                         sys__mgr7__ready               ;
  input                                         sys__mgr7__complete            ;
  // General control and status                                                   
  output                                        mgr8__sys__allSynchronized     ;
  input                                         sys__mgr8__thisSynchronized    ;
  input                                         sys__mgr8__ready               ;
  input                                         sys__mgr8__complete            ;
  // General control and status                                                   
  output                                        mgr9__sys__allSynchronized     ;
  input                                         sys__mgr9__thisSynchronized    ;
  input                                         sys__mgr9__ready               ;
  input                                         sys__mgr9__complete            ;
  // General control and status                                                   
  output                                        mgr10__sys__allSynchronized     ;
  input                                         sys__mgr10__thisSynchronized    ;
  input                                         sys__mgr10__ready               ;
  input                                         sys__mgr10__complete            ;
  // General control and status                                                   
  output                                        mgr11__sys__allSynchronized     ;
  input                                         sys__mgr11__thisSynchronized    ;
  input                                         sys__mgr11__ready               ;
  input                                         sys__mgr11__complete            ;
  // General control and status                                                   
  output                                        mgr12__sys__allSynchronized     ;
  input                                         sys__mgr12__thisSynchronized    ;
  input                                         sys__mgr12__ready               ;
  input                                         sys__mgr12__complete            ;
  // General control and status                                                   
  output                                        mgr13__sys__allSynchronized     ;
  input                                         sys__mgr13__thisSynchronized    ;
  input                                         sys__mgr13__ready               ;
  input                                         sys__mgr13__complete            ;
  // General control and status                                                   
  output                                        mgr14__sys__allSynchronized     ;
  input                                         sys__mgr14__thisSynchronized    ;
  input                                         sys__mgr14__ready               ;
  input                                         sys__mgr14__complete            ;
  // General control and status                                                   
  output                                        mgr15__sys__allSynchronized     ;
  input                                         sys__mgr15__thisSynchronized    ;
  input                                         sys__mgr15__ready               ;
  input                                         sys__mgr15__complete            ;
  // General control and status                                                   
  output                                        mgr16__sys__allSynchronized     ;
  input                                         sys__mgr16__thisSynchronized    ;
  input                                         sys__mgr16__ready               ;
  input                                         sys__mgr16__complete            ;
  // General control and status                                                   
  output                                        mgr17__sys__allSynchronized     ;
  input                                         sys__mgr17__thisSynchronized    ;
  input                                         sys__mgr17__ready               ;
  input                                         sys__mgr17__complete            ;
  // General control and status                                                   
  output                                        mgr18__sys__allSynchronized     ;
  input                                         sys__mgr18__thisSynchronized    ;
  input                                         sys__mgr18__ready               ;
  input                                         sys__mgr18__complete            ;
  // General control and status                                                   
  output                                        mgr19__sys__allSynchronized     ;
  input                                         sys__mgr19__thisSynchronized    ;
  input                                         sys__mgr19__ready               ;
  input                                         sys__mgr19__complete            ;
  // General control and status                                                   
  output                                        mgr20__sys__allSynchronized     ;
  input                                         sys__mgr20__thisSynchronized    ;
  input                                         sys__mgr20__ready               ;
  input                                         sys__mgr20__complete            ;
  // General control and status                                                   
  output                                        mgr21__sys__allSynchronized     ;
  input                                         sys__mgr21__thisSynchronized    ;
  input                                         sys__mgr21__ready               ;
  input                                         sys__mgr21__complete            ;
  // General control and status                                                   
  output                                        mgr22__sys__allSynchronized     ;
  input                                         sys__mgr22__thisSynchronized    ;
  input                                         sys__mgr22__ready               ;
  input                                         sys__mgr22__complete            ;
  // General control and status                                                   
  output                                        mgr23__sys__allSynchronized     ;
  input                                         sys__mgr23__thisSynchronized    ;
  input                                         sys__mgr23__ready               ;
  input                                         sys__mgr23__complete            ;
  // General control and status                                                   
  output                                        mgr24__sys__allSynchronized     ;
  input                                         sys__mgr24__thisSynchronized    ;
  input                                         sys__mgr24__ready               ;
  input                                         sys__mgr24__complete            ;
  // General control and status                                                   
  output                                        mgr25__sys__allSynchronized     ;
  input                                         sys__mgr25__thisSynchronized    ;
  input                                         sys__mgr25__ready               ;
  input                                         sys__mgr25__complete            ;
  // General control and status                                                   
  output                                        mgr26__sys__allSynchronized     ;
  input                                         sys__mgr26__thisSynchronized    ;
  input                                         sys__mgr26__ready               ;
  input                                         sys__mgr26__complete            ;
  // General control and status                                                   
  output                                        mgr27__sys__allSynchronized     ;
  input                                         sys__mgr27__thisSynchronized    ;
  input                                         sys__mgr27__ready               ;
  input                                         sys__mgr27__complete            ;
  // General control and status                                                   
  output                                        mgr28__sys__allSynchronized     ;
  input                                         sys__mgr28__thisSynchronized    ;
  input                                         sys__mgr28__ready               ;
  input                                         sys__mgr28__complete            ;
  // General control and status                                                   
  output                                        mgr29__sys__allSynchronized     ;
  input                                         sys__mgr29__thisSynchronized    ;
  input                                         sys__mgr29__ready               ;
  input                                         sys__mgr29__complete            ;
  // General control and status                                                   
  output                                        mgr30__sys__allSynchronized     ;
  input                                         sys__mgr30__thisSynchronized    ;
  input                                         sys__mgr30__ready               ;
  input                                         sys__mgr30__complete            ;
  // General control and status                                                   
  output                                        mgr31__sys__allSynchronized     ;
  input                                         sys__mgr31__thisSynchronized    ;
  input                                         sys__mgr31__ready               ;
  input                                         sys__mgr31__complete            ;
  // General control and status                                                   
  output                                        mgr32__sys__allSynchronized     ;
  input                                         sys__mgr32__thisSynchronized    ;
  input                                         sys__mgr32__ready               ;
  input                                         sys__mgr32__complete            ;
  // General control and status                                                   
  output                                        mgr33__sys__allSynchronized     ;
  input                                         sys__mgr33__thisSynchronized    ;
  input                                         sys__mgr33__ready               ;
  input                                         sys__mgr33__complete            ;
  // General control and status                                                   
  output                                        mgr34__sys__allSynchronized     ;
  input                                         sys__mgr34__thisSynchronized    ;
  input                                         sys__mgr34__ready               ;
  input                                         sys__mgr34__complete            ;
  // General control and status                                                   
  output                                        mgr35__sys__allSynchronized     ;
  input                                         sys__mgr35__thisSynchronized    ;
  input                                         sys__mgr35__ready               ;
  input                                         sys__mgr35__complete            ;
  // General control and status                                                   
  output                                        mgr36__sys__allSynchronized     ;
  input                                         sys__mgr36__thisSynchronized    ;
  input                                         sys__mgr36__ready               ;
  input                                         sys__mgr36__complete            ;
  // General control and status                                                   
  output                                        mgr37__sys__allSynchronized     ;
  input                                         sys__mgr37__thisSynchronized    ;
  input                                         sys__mgr37__ready               ;
  input                                         sys__mgr37__complete            ;
  // General control and status                                                   
  output                                        mgr38__sys__allSynchronized     ;
  input                                         sys__mgr38__thisSynchronized    ;
  input                                         sys__mgr38__ready               ;
  input                                         sys__mgr38__complete            ;
  // General control and status                                                   
  output                                        mgr39__sys__allSynchronized     ;
  input                                         sys__mgr39__thisSynchronized    ;
  input                                         sys__mgr39__ready               ;
  input                                         sys__mgr39__complete            ;
  // General control and status                                                   
  output                                        mgr40__sys__allSynchronized     ;
  input                                         sys__mgr40__thisSynchronized    ;
  input                                         sys__mgr40__ready               ;
  input                                         sys__mgr40__complete            ;
  // General control and status                                                   
  output                                        mgr41__sys__allSynchronized     ;
  input                                         sys__mgr41__thisSynchronized    ;
  input                                         sys__mgr41__ready               ;
  input                                         sys__mgr41__complete            ;
  // General control and status                                                   
  output                                        mgr42__sys__allSynchronized     ;
  input                                         sys__mgr42__thisSynchronized    ;
  input                                         sys__mgr42__ready               ;
  input                                         sys__mgr42__complete            ;
  // General control and status                                                   
  output                                        mgr43__sys__allSynchronized     ;
  input                                         sys__mgr43__thisSynchronized    ;
  input                                         sys__mgr43__ready               ;
  input                                         sys__mgr43__complete            ;
  // General control and status                                                   
  output                                        mgr44__sys__allSynchronized     ;
  input                                         sys__mgr44__thisSynchronized    ;
  input                                         sys__mgr44__ready               ;
  input                                         sys__mgr44__complete            ;
  // General control and status                                                   
  output                                        mgr45__sys__allSynchronized     ;
  input                                         sys__mgr45__thisSynchronized    ;
  input                                         sys__mgr45__ready               ;
  input                                         sys__mgr45__complete            ;
  // General control and status                                                   
  output                                        mgr46__sys__allSynchronized     ;
  input                                         sys__mgr46__thisSynchronized    ;
  input                                         sys__mgr46__ready               ;
  input                                         sys__mgr46__complete            ;
  // General control and status                                                   
  output                                        mgr47__sys__allSynchronized     ;
  input                                         sys__mgr47__thisSynchronized    ;
  input                                         sys__mgr47__ready               ;
  input                                         sys__mgr47__complete            ;
  // General control and status                                                   
  output                                        mgr48__sys__allSynchronized     ;
  input                                         sys__mgr48__thisSynchronized    ;
  input                                         sys__mgr48__ready               ;
  input                                         sys__mgr48__complete            ;
  // General control and status                                                   
  output                                        mgr49__sys__allSynchronized     ;
  input                                         sys__mgr49__thisSynchronized    ;
  input                                         sys__mgr49__ready               ;
  input                                         sys__mgr49__complete            ;
  // General control and status                                                   
  output                                        mgr50__sys__allSynchronized     ;
  input                                         sys__mgr50__thisSynchronized    ;
  input                                         sys__mgr50__ready               ;
  input                                         sys__mgr50__complete            ;
  // General control and status                                                   
  output                                        mgr51__sys__allSynchronized     ;
  input                                         sys__mgr51__thisSynchronized    ;
  input                                         sys__mgr51__ready               ;
  input                                         sys__mgr51__complete            ;
  // General control and status                                                   
  output                                        mgr52__sys__allSynchronized     ;
  input                                         sys__mgr52__thisSynchronized    ;
  input                                         sys__mgr52__ready               ;
  input                                         sys__mgr52__complete            ;
  // General control and status                                                   
  output                                        mgr53__sys__allSynchronized     ;
  input                                         sys__mgr53__thisSynchronized    ;
  input                                         sys__mgr53__ready               ;
  input                                         sys__mgr53__complete            ;
  // General control and status                                                   
  output                                        mgr54__sys__allSynchronized     ;
  input                                         sys__mgr54__thisSynchronized    ;
  input                                         sys__mgr54__ready               ;
  input                                         sys__mgr54__complete            ;
  // General control and status                                                   
  output                                        mgr55__sys__allSynchronized     ;
  input                                         sys__mgr55__thisSynchronized    ;
  input                                         sys__mgr55__ready               ;
  input                                         sys__mgr55__complete            ;
  // General control and status                                                   
  output                                        mgr56__sys__allSynchronized     ;
  input                                         sys__mgr56__thisSynchronized    ;
  input                                         sys__mgr56__ready               ;
  input                                         sys__mgr56__complete            ;
  // General control and status                                                   
  output                                        mgr57__sys__allSynchronized     ;
  input                                         sys__mgr57__thisSynchronized    ;
  input                                         sys__mgr57__ready               ;
  input                                         sys__mgr57__complete            ;
  // General control and status                                                   
  output                                        mgr58__sys__allSynchronized     ;
  input                                         sys__mgr58__thisSynchronized    ;
  input                                         sys__mgr58__ready               ;
  input                                         sys__mgr58__complete            ;
  // General control and status                                                   
  output                                        mgr59__sys__allSynchronized     ;
  input                                         sys__mgr59__thisSynchronized    ;
  input                                         sys__mgr59__ready               ;
  input                                         sys__mgr59__complete            ;
  // General control and status                                                   
  output                                        mgr60__sys__allSynchronized     ;
  input                                         sys__mgr60__thisSynchronized    ;
  input                                         sys__mgr60__ready               ;
  input                                         sys__mgr60__complete            ;
  // General control and status                                                   
  output                                        mgr61__sys__allSynchronized     ;
  input                                         sys__mgr61__thisSynchronized    ;
  input                                         sys__mgr61__ready               ;
  input                                         sys__mgr61__complete            ;
  // General control and status                                                   
  output                                        mgr62__sys__allSynchronized     ;
  input                                         sys__mgr62__thisSynchronized    ;
  input                                         sys__mgr62__ready               ;
  input                                         sys__mgr62__complete            ;
  // General control and status                                                   
  output                                        mgr63__sys__allSynchronized     ;
  input                                         sys__mgr63__thisSynchronized    ;
  input                                         sys__mgr63__ready               ;
  input                                         sys__mgr63__complete            ;