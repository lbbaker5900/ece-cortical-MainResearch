
            // General control and status                  
            sys__pe0__allSynchronized                    ,
            pe0__sys__thisSynchronized                   ,
            pe0__sys__ready                              ,
            pe0__sys__complete                           ,
            // General control and status                  
            sys__pe1__allSynchronized                    ,
            pe1__sys__thisSynchronized                   ,
            pe1__sys__ready                              ,
            pe1__sys__complete                           ,
            // General control and status                  
            sys__pe2__allSynchronized                    ,
            pe2__sys__thisSynchronized                   ,
            pe2__sys__ready                              ,
            pe2__sys__complete                           ,
            // General control and status                  
            sys__pe3__allSynchronized                    ,
            pe3__sys__thisSynchronized                   ,
            pe3__sys__ready                              ,
            pe3__sys__complete                           ,