
    // MGR0, Port0 next hop mask                 
    assign mgr_inst[0].sys__mgr__port_destinationMask [0]    = `MGR_NOC_CONT_MGR0_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR0, Port1 next hop mask                 
    assign mgr_inst[0].sys__mgr__port_destinationMask [1]    = `MGR_NOC_CONT_MGR0_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR0, Port2 next hop mask                 
    assign mgr_inst[0].sys__mgr__port_destinationMask [2]    = `MGR_NOC_CONT_MGR0_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR0, Port3 next hop mask                 
    assign mgr_inst[0].sys__mgr__port_destinationMask [3]    = `MGR_NOC_CONT_MGR0_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR1, Port0 next hop mask                 
    assign mgr_inst[1].sys__mgr__port_destinationMask [0]    = `MGR_NOC_CONT_MGR1_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR1, Port1 next hop mask                 
    assign mgr_inst[1].sys__mgr__port_destinationMask [1]    = `MGR_NOC_CONT_MGR1_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR1, Port2 next hop mask                 
    assign mgr_inst[1].sys__mgr__port_destinationMask [2]    = `MGR_NOC_CONT_MGR1_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR1, Port3 next hop mask                 
    assign mgr_inst[1].sys__mgr__port_destinationMask [3]    = `MGR_NOC_CONT_MGR1_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR2, Port0 next hop mask                 
    assign mgr_inst[2].sys__mgr__port_destinationMask [0]    = `MGR_NOC_CONT_MGR2_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR2, Port1 next hop mask                 
    assign mgr_inst[2].sys__mgr__port_destinationMask [1]    = `MGR_NOC_CONT_MGR2_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR2, Port2 next hop mask                 
    assign mgr_inst[2].sys__mgr__port_destinationMask [2]    = `MGR_NOC_CONT_MGR2_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR2, Port3 next hop mask                 
    assign mgr_inst[2].sys__mgr__port_destinationMask [3]    = `MGR_NOC_CONT_MGR2_PORT3_DESTINATION_MGR_BITMASK ;
    // MGR3, Port0 next hop mask                 
    assign mgr_inst[3].sys__mgr__port_destinationMask [0]    = `MGR_NOC_CONT_MGR3_PORT0_DESTINATION_MGR_BITMASK ;
    // MGR3, Port1 next hop mask                 
    assign mgr_inst[3].sys__mgr__port_destinationMask [1]    = `MGR_NOC_CONT_MGR3_PORT1_DESTINATION_MGR_BITMASK ;
    // MGR3, Port2 next hop mask                 
    assign mgr_inst[3].sys__mgr__port_destinationMask [2]    = `MGR_NOC_CONT_MGR3_PORT2_DESTINATION_MGR_BITMASK ;
    // MGR3, Port3 next hop mask                 
    assign mgr_inst[3].sys__mgr__port_destinationMask [3]    = `MGR_NOC_CONT_MGR3_PORT3_DESTINATION_MGR_BITMASK ;