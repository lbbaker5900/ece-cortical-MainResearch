
    output                                         stu__mgr0__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr0__cntl           ;
    input                                          mgr0__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr0__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr0__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr0__oob_data       ;

    input                                          pe0__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe0__stu__cntl           ;
    output                                         stu__pe0__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe0__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe0__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe0__stu__oob_data       ;

    output                                         stu__mgr1__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr1__cntl           ;
    input                                          mgr1__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr1__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr1__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr1__oob_data       ;

    input                                          pe1__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe1__stu__cntl           ;
    output                                         stu__pe1__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe1__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe1__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe1__stu__oob_data       ;

    output                                         stu__mgr2__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr2__cntl           ;
    input                                          mgr2__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr2__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr2__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr2__oob_data       ;

    input                                          pe2__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe2__stu__cntl           ;
    output                                         stu__pe2__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe2__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe2__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe2__stu__oob_data       ;

    output                                         stu__mgr3__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr3__cntl           ;
    input                                          mgr3__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr3__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr3__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr3__oob_data       ;

    input                                          pe3__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe3__stu__cntl           ;
    output                                         stu__pe3__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe3__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe3__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe3__stu__oob_data       ;

    output                                         stu__mgr4__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr4__cntl           ;
    input                                          mgr4__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr4__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr4__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr4__oob_data       ;

    input                                          pe4__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe4__stu__cntl           ;
    output                                         stu__pe4__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe4__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe4__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe4__stu__oob_data       ;

    output                                         stu__mgr5__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr5__cntl           ;
    input                                          mgr5__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr5__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr5__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr5__oob_data       ;

    input                                          pe5__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe5__stu__cntl           ;
    output                                         stu__pe5__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe5__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe5__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe5__stu__oob_data       ;

    output                                         stu__mgr6__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr6__cntl           ;
    input                                          mgr6__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr6__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr6__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr6__oob_data       ;

    input                                          pe6__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe6__stu__cntl           ;
    output                                         stu__pe6__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe6__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe6__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe6__stu__oob_data       ;

    output                                         stu__mgr7__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr7__cntl           ;
    input                                          mgr7__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr7__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr7__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr7__oob_data       ;

    input                                          pe7__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe7__stu__cntl           ;
    output                                         stu__pe7__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe7__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe7__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe7__stu__oob_data       ;

    output                                         stu__mgr8__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr8__cntl           ;
    input                                          mgr8__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr8__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr8__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr8__oob_data       ;

    input                                          pe8__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe8__stu__cntl           ;
    output                                         stu__pe8__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe8__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe8__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe8__stu__oob_data       ;

    output                                         stu__mgr9__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr9__cntl           ;
    input                                          mgr9__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr9__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr9__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr9__oob_data       ;

    input                                          pe9__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe9__stu__cntl           ;
    output                                         stu__pe9__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe9__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe9__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe9__stu__oob_data       ;

    output                                         stu__mgr10__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr10__cntl           ;
    input                                          mgr10__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr10__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr10__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr10__oob_data       ;

    input                                          pe10__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe10__stu__cntl           ;
    output                                         stu__pe10__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe10__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe10__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe10__stu__oob_data       ;

    output                                         stu__mgr11__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr11__cntl           ;
    input                                          mgr11__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr11__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr11__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr11__oob_data       ;

    input                                          pe11__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe11__stu__cntl           ;
    output                                         stu__pe11__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe11__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe11__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe11__stu__oob_data       ;

    output                                         stu__mgr12__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr12__cntl           ;
    input                                          mgr12__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr12__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr12__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr12__oob_data       ;

    input                                          pe12__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe12__stu__cntl           ;
    output                                         stu__pe12__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe12__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe12__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe12__stu__oob_data       ;

    output                                         stu__mgr13__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr13__cntl           ;
    input                                          mgr13__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr13__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr13__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr13__oob_data       ;

    input                                          pe13__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe13__stu__cntl           ;
    output                                         stu__pe13__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe13__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe13__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe13__stu__oob_data       ;

    output                                         stu__mgr14__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr14__cntl           ;
    input                                          mgr14__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr14__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr14__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr14__oob_data       ;

    input                                          pe14__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe14__stu__cntl           ;
    output                                         stu__pe14__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe14__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe14__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe14__stu__oob_data       ;

    output                                         stu__mgr15__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr15__cntl           ;
    input                                          mgr15__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr15__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr15__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr15__oob_data       ;

    input                                          pe15__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe15__stu__cntl           ;
    output                                         stu__pe15__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe15__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe15__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe15__stu__oob_data       ;

    output                                         stu__mgr16__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr16__cntl           ;
    input                                          mgr16__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr16__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr16__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr16__oob_data       ;

    input                                          pe16__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe16__stu__cntl           ;
    output                                         stu__pe16__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe16__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe16__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe16__stu__oob_data       ;

    output                                         stu__mgr17__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr17__cntl           ;
    input                                          mgr17__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr17__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr17__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr17__oob_data       ;

    input                                          pe17__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe17__stu__cntl           ;
    output                                         stu__pe17__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe17__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe17__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe17__stu__oob_data       ;

    output                                         stu__mgr18__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr18__cntl           ;
    input                                          mgr18__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr18__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr18__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr18__oob_data       ;

    input                                          pe18__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe18__stu__cntl           ;
    output                                         stu__pe18__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe18__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe18__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe18__stu__oob_data       ;

    output                                         stu__mgr19__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr19__cntl           ;
    input                                          mgr19__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr19__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr19__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr19__oob_data       ;

    input                                          pe19__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe19__stu__cntl           ;
    output                                         stu__pe19__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe19__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe19__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe19__stu__oob_data       ;

    output                                         stu__mgr20__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr20__cntl           ;
    input                                          mgr20__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr20__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr20__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr20__oob_data       ;

    input                                          pe20__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe20__stu__cntl           ;
    output                                         stu__pe20__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe20__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe20__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe20__stu__oob_data       ;

    output                                         stu__mgr21__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr21__cntl           ;
    input                                          mgr21__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr21__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr21__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr21__oob_data       ;

    input                                          pe21__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe21__stu__cntl           ;
    output                                         stu__pe21__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe21__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe21__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe21__stu__oob_data       ;

    output                                         stu__mgr22__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr22__cntl           ;
    input                                          mgr22__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr22__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr22__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr22__oob_data       ;

    input                                          pe22__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe22__stu__cntl           ;
    output                                         stu__pe22__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe22__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe22__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe22__stu__oob_data       ;

    output                                         stu__mgr23__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr23__cntl           ;
    input                                          mgr23__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr23__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr23__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr23__oob_data       ;

    input                                          pe23__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe23__stu__cntl           ;
    output                                         stu__pe23__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe23__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe23__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe23__stu__oob_data       ;

    output                                         stu__mgr24__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr24__cntl           ;
    input                                          mgr24__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr24__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr24__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr24__oob_data       ;

    input                                          pe24__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe24__stu__cntl           ;
    output                                         stu__pe24__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe24__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe24__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe24__stu__oob_data       ;

    output                                         stu__mgr25__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr25__cntl           ;
    input                                          mgr25__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr25__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr25__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr25__oob_data       ;

    input                                          pe25__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe25__stu__cntl           ;
    output                                         stu__pe25__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe25__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe25__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe25__stu__oob_data       ;

    output                                         stu__mgr26__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr26__cntl           ;
    input                                          mgr26__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr26__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr26__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr26__oob_data       ;

    input                                          pe26__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe26__stu__cntl           ;
    output                                         stu__pe26__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe26__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe26__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe26__stu__oob_data       ;

    output                                         stu__mgr27__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr27__cntl           ;
    input                                          mgr27__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr27__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr27__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr27__oob_data       ;

    input                                          pe27__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe27__stu__cntl           ;
    output                                         stu__pe27__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe27__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe27__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe27__stu__oob_data       ;

    output                                         stu__mgr28__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr28__cntl           ;
    input                                          mgr28__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr28__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr28__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr28__oob_data       ;

    input                                          pe28__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe28__stu__cntl           ;
    output                                         stu__pe28__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe28__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe28__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe28__stu__oob_data       ;

    output                                         stu__mgr29__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr29__cntl           ;
    input                                          mgr29__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr29__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr29__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr29__oob_data       ;

    input                                          pe29__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe29__stu__cntl           ;
    output                                         stu__pe29__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe29__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe29__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe29__stu__oob_data       ;

    output                                         stu__mgr30__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr30__cntl           ;
    input                                          mgr30__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr30__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr30__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr30__oob_data       ;

    input                                          pe30__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe30__stu__cntl           ;
    output                                         stu__pe30__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe30__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe30__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe30__stu__oob_data       ;

    output                                         stu__mgr31__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr31__cntl           ;
    input                                          mgr31__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr31__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr31__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr31__oob_data       ;

    input                                          pe31__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe31__stu__cntl           ;
    output                                         stu__pe31__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe31__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe31__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe31__stu__oob_data       ;

    output                                         stu__mgr32__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr32__cntl           ;
    input                                          mgr32__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr32__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr32__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr32__oob_data       ;

    input                                          pe32__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe32__stu__cntl           ;
    output                                         stu__pe32__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe32__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe32__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe32__stu__oob_data       ;

    output                                         stu__mgr33__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr33__cntl           ;
    input                                          mgr33__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr33__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr33__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr33__oob_data       ;

    input                                          pe33__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe33__stu__cntl           ;
    output                                         stu__pe33__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe33__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe33__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe33__stu__oob_data       ;

    output                                         stu__mgr34__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr34__cntl           ;
    input                                          mgr34__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr34__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr34__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr34__oob_data       ;

    input                                          pe34__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe34__stu__cntl           ;
    output                                         stu__pe34__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe34__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe34__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe34__stu__oob_data       ;

    output                                         stu__mgr35__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr35__cntl           ;
    input                                          mgr35__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr35__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr35__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr35__oob_data       ;

    input                                          pe35__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe35__stu__cntl           ;
    output                                         stu__pe35__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe35__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe35__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe35__stu__oob_data       ;

    output                                         stu__mgr36__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr36__cntl           ;
    input                                          mgr36__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr36__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr36__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr36__oob_data       ;

    input                                          pe36__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe36__stu__cntl           ;
    output                                         stu__pe36__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe36__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe36__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe36__stu__oob_data       ;

    output                                         stu__mgr37__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr37__cntl           ;
    input                                          mgr37__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr37__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr37__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr37__oob_data       ;

    input                                          pe37__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe37__stu__cntl           ;
    output                                         stu__pe37__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe37__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe37__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe37__stu__oob_data       ;

    output                                         stu__mgr38__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr38__cntl           ;
    input                                          mgr38__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr38__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr38__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr38__oob_data       ;

    input                                          pe38__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe38__stu__cntl           ;
    output                                         stu__pe38__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe38__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe38__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe38__stu__oob_data       ;

    output                                         stu__mgr39__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr39__cntl           ;
    input                                          mgr39__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr39__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr39__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr39__oob_data       ;

    input                                          pe39__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe39__stu__cntl           ;
    output                                         stu__pe39__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe39__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe39__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe39__stu__oob_data       ;

    output                                         stu__mgr40__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr40__cntl           ;
    input                                          mgr40__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr40__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr40__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr40__oob_data       ;

    input                                          pe40__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe40__stu__cntl           ;
    output                                         stu__pe40__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe40__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe40__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe40__stu__oob_data       ;

    output                                         stu__mgr41__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr41__cntl           ;
    input                                          mgr41__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr41__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr41__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr41__oob_data       ;

    input                                          pe41__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe41__stu__cntl           ;
    output                                         stu__pe41__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe41__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe41__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe41__stu__oob_data       ;

    output                                         stu__mgr42__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr42__cntl           ;
    input                                          mgr42__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr42__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr42__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr42__oob_data       ;

    input                                          pe42__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe42__stu__cntl           ;
    output                                         stu__pe42__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe42__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe42__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe42__stu__oob_data       ;

    output                                         stu__mgr43__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr43__cntl           ;
    input                                          mgr43__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr43__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr43__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr43__oob_data       ;

    input                                          pe43__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe43__stu__cntl           ;
    output                                         stu__pe43__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe43__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe43__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe43__stu__oob_data       ;

    output                                         stu__mgr44__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr44__cntl           ;
    input                                          mgr44__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr44__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr44__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr44__oob_data       ;

    input                                          pe44__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe44__stu__cntl           ;
    output                                         stu__pe44__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe44__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe44__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe44__stu__oob_data       ;

    output                                         stu__mgr45__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr45__cntl           ;
    input                                          mgr45__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr45__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr45__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr45__oob_data       ;

    input                                          pe45__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe45__stu__cntl           ;
    output                                         stu__pe45__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe45__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe45__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe45__stu__oob_data       ;

    output                                         stu__mgr46__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr46__cntl           ;
    input                                          mgr46__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr46__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr46__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr46__oob_data       ;

    input                                          pe46__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe46__stu__cntl           ;
    output                                         stu__pe46__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe46__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe46__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe46__stu__oob_data       ;

    output                                         stu__mgr47__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr47__cntl           ;
    input                                          mgr47__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr47__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr47__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr47__oob_data       ;

    input                                          pe47__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe47__stu__cntl           ;
    output                                         stu__pe47__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe47__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe47__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe47__stu__oob_data       ;

    output                                         stu__mgr48__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr48__cntl           ;
    input                                          mgr48__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr48__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr48__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr48__oob_data       ;

    input                                          pe48__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe48__stu__cntl           ;
    output                                         stu__pe48__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe48__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe48__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe48__stu__oob_data       ;

    output                                         stu__mgr49__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr49__cntl           ;
    input                                          mgr49__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr49__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr49__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr49__oob_data       ;

    input                                          pe49__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe49__stu__cntl           ;
    output                                         stu__pe49__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe49__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe49__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe49__stu__oob_data       ;

    output                                         stu__mgr50__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr50__cntl           ;
    input                                          mgr50__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr50__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr50__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr50__oob_data       ;

    input                                          pe50__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe50__stu__cntl           ;
    output                                         stu__pe50__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe50__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe50__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe50__stu__oob_data       ;

    output                                         stu__mgr51__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr51__cntl           ;
    input                                          mgr51__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr51__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr51__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr51__oob_data       ;

    input                                          pe51__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe51__stu__cntl           ;
    output                                         stu__pe51__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe51__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe51__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe51__stu__oob_data       ;

    output                                         stu__mgr52__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr52__cntl           ;
    input                                          mgr52__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr52__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr52__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr52__oob_data       ;

    input                                          pe52__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe52__stu__cntl           ;
    output                                         stu__pe52__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe52__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe52__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe52__stu__oob_data       ;

    output                                         stu__mgr53__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr53__cntl           ;
    input                                          mgr53__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr53__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr53__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr53__oob_data       ;

    input                                          pe53__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe53__stu__cntl           ;
    output                                         stu__pe53__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe53__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe53__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe53__stu__oob_data       ;

    output                                         stu__mgr54__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr54__cntl           ;
    input                                          mgr54__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr54__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr54__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr54__oob_data       ;

    input                                          pe54__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe54__stu__cntl           ;
    output                                         stu__pe54__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe54__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe54__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe54__stu__oob_data       ;

    output                                         stu__mgr55__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr55__cntl           ;
    input                                          mgr55__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr55__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr55__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr55__oob_data       ;

    input                                          pe55__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe55__stu__cntl           ;
    output                                         stu__pe55__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe55__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe55__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe55__stu__oob_data       ;

    output                                         stu__mgr56__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr56__cntl           ;
    input                                          mgr56__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr56__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr56__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr56__oob_data       ;

    input                                          pe56__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe56__stu__cntl           ;
    output                                         stu__pe56__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe56__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe56__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe56__stu__oob_data       ;

    output                                         stu__mgr57__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr57__cntl           ;
    input                                          mgr57__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr57__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr57__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr57__oob_data       ;

    input                                          pe57__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe57__stu__cntl           ;
    output                                         stu__pe57__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe57__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe57__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe57__stu__oob_data       ;

    output                                         stu__mgr58__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr58__cntl           ;
    input                                          mgr58__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr58__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr58__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr58__oob_data       ;

    input                                          pe58__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe58__stu__cntl           ;
    output                                         stu__pe58__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe58__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe58__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe58__stu__oob_data       ;

    output                                         stu__mgr59__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr59__cntl           ;
    input                                          mgr59__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr59__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr59__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr59__oob_data       ;

    input                                          pe59__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe59__stu__cntl           ;
    output                                         stu__pe59__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe59__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe59__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe59__stu__oob_data       ;

    output                                         stu__mgr60__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr60__cntl           ;
    input                                          mgr60__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr60__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr60__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr60__oob_data       ;

    input                                          pe60__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe60__stu__cntl           ;
    output                                         stu__pe60__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe60__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe60__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe60__stu__oob_data       ;

    output                                         stu__mgr61__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr61__cntl           ;
    input                                          mgr61__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr61__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr61__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr61__oob_data       ;

    input                                          pe61__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe61__stu__cntl           ;
    output                                         stu__pe61__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe61__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe61__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe61__stu__oob_data       ;

    output                                         stu__mgr62__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr62__cntl           ;
    input                                          mgr62__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr62__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr62__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr62__oob_data       ;

    input                                          pe62__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe62__stu__cntl           ;
    output                                         stu__pe62__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe62__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe62__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe62__stu__oob_data       ;

    output                                         stu__mgr63__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr63__cntl           ;
    input                                          mgr63__stu__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr63__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr63__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr63__oob_data       ;

    input                                          pe63__stu__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       pe63__stu__cntl           ;
    output                                         stu__pe63__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       pe63__stu__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       pe63__stu__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe63__stu__oob_data       ;

