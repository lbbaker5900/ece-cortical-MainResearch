
  input                                    reg__scntl__lane0_ready    ;
  output                                   scntl__reg__lane0_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane0_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane0_data     ;

  input                                    reg__scntl__lane1_ready    ;
  output                                   scntl__reg__lane1_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane1_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane1_data     ;

  input                                    reg__scntl__lane2_ready    ;
  output                                   scntl__reg__lane2_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane2_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane2_data     ;

  input                                    reg__scntl__lane3_ready    ;
  output                                   scntl__reg__lane3_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane3_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane3_data     ;

  input                                    reg__scntl__lane4_ready    ;
  output                                   scntl__reg__lane4_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane4_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane4_data     ;

  input                                    reg__scntl__lane5_ready    ;
  output                                   scntl__reg__lane5_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane5_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane5_data     ;

  input                                    reg__scntl__lane6_ready    ;
  output                                   scntl__reg__lane6_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane6_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane6_data     ;

  input                                    reg__scntl__lane7_ready    ;
  output                                   scntl__reg__lane7_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane7_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane7_data     ;

  input                                    reg__scntl__lane8_ready    ;
  output                                   scntl__reg__lane8_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane8_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane8_data     ;

  input                                    reg__scntl__lane9_ready    ;
  output                                   scntl__reg__lane9_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane9_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane9_data     ;

  input                                    reg__scntl__lane10_ready    ;
  output                                   scntl__reg__lane10_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane10_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane10_data     ;

  input                                    reg__scntl__lane11_ready    ;
  output                                   scntl__reg__lane11_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane11_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane11_data     ;

  input                                    reg__scntl__lane12_ready    ;
  output                                   scntl__reg__lane12_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane12_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane12_data     ;

  input                                    reg__scntl__lane13_ready    ;
  output                                   scntl__reg__lane13_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane13_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane13_data     ;

  input                                    reg__scntl__lane14_ready    ;
  output                                   scntl__reg__lane14_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane14_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane14_data     ;

  input                                    reg__scntl__lane15_ready    ;
  output                                   scntl__reg__lane15_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane15_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane15_data     ;

  input                                    reg__scntl__lane16_ready    ;
  output                                   scntl__reg__lane16_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane16_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane16_data     ;

  input                                    reg__scntl__lane17_ready    ;
  output                                   scntl__reg__lane17_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane17_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane17_data     ;

  input                                    reg__scntl__lane18_ready    ;
  output                                   scntl__reg__lane18_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane18_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane18_data     ;

  input                                    reg__scntl__lane19_ready    ;
  output                                   scntl__reg__lane19_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane19_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane19_data     ;

  input                                    reg__scntl__lane20_ready    ;
  output                                   scntl__reg__lane20_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane20_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane20_data     ;

  input                                    reg__scntl__lane21_ready    ;
  output                                   scntl__reg__lane21_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane21_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane21_data     ;

  input                                    reg__scntl__lane22_ready    ;
  output                                   scntl__reg__lane22_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane22_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane22_data     ;

  input                                    reg__scntl__lane23_ready    ;
  output                                   scntl__reg__lane23_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane23_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane23_data     ;

  input                                    reg__scntl__lane24_ready    ;
  output                                   scntl__reg__lane24_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane24_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane24_data     ;

  input                                    reg__scntl__lane25_ready    ;
  output                                   scntl__reg__lane25_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane25_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane25_data     ;

  input                                    reg__scntl__lane26_ready    ;
  output                                   scntl__reg__lane26_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane26_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane26_data     ;

  input                                    reg__scntl__lane27_ready    ;
  output                                   scntl__reg__lane27_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane27_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane27_data     ;

  input                                    reg__scntl__lane28_ready    ;
  output                                   scntl__reg__lane28_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane28_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane28_data     ;

  input                                    reg__scntl__lane29_ready    ;
  output                                   scntl__reg__lane29_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane29_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane29_data     ;

  input                                    reg__scntl__lane30_ready    ;
  output                                   scntl__reg__lane30_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane30_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane30_data     ;

  input                                    reg__scntl__lane31_ready    ;
  output                                   scntl__reg__lane31_valid    ;
  output  [`COMMON_STD_INTF_CNTL_RANGE  ]  scntl__reg__lane31_cntl     ;
  output  [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane31_data     ;

