
  // NoC port 0
  reg                                      pe__noc__port0_valid           ;
  wire   [`COMMON_STD_INTF_CNTL_RANGE ]  pe__noc__port0_cntl            ;
  wire   [`NOC_CONT_NOC_PORT_DATA_RANGE ]  pe__noc__port0_data            ;
  wire                                     noc__pe__port0_fc              ;
  wire                                     noc__pe__port0_valid           ;
  wire   [`COMMON_STD_INTF_CNTL_RANGE ]  noc__pe__port0_cntl            ;
  wire   [`NOC_CONT_NOC_PORT_DATA_RANGE ]  noc__pe__port0_data            ;
  wire                                     pe__noc__port0_fc              ;
  wire   [`PE_PE_ID_BITMASK_RANGE       ]  sys__pe__port0_destinationMask ;

  // NoC port 1
  reg                                      pe__noc__port1_valid           ;
  wire   [`COMMON_STD_INTF_CNTL_RANGE ]  pe__noc__port1_cntl            ;
  wire   [`NOC_CONT_NOC_PORT_DATA_RANGE ]  pe__noc__port1_data            ;
  wire                                     noc__pe__port1_fc              ;
  wire                                     noc__pe__port1_valid           ;
  wire   [`COMMON_STD_INTF_CNTL_RANGE ]  noc__pe__port1_cntl            ;
  wire   [`NOC_CONT_NOC_PORT_DATA_RANGE ]  noc__pe__port1_data            ;
  wire                                     pe__noc__port1_fc              ;
  wire   [`PE_PE_ID_BITMASK_RANGE       ]  sys__pe__port1_destinationMask ;

  // NoC port 2
  reg                                      pe__noc__port2_valid           ;
  wire   [`COMMON_STD_INTF_CNTL_RANGE ]  pe__noc__port2_cntl            ;
  wire   [`NOC_CONT_NOC_PORT_DATA_RANGE ]  pe__noc__port2_data            ;
  wire                                     noc__pe__port2_fc              ;
  wire                                     noc__pe__port2_valid           ;
  wire   [`COMMON_STD_INTF_CNTL_RANGE ]  noc__pe__port2_cntl            ;
  wire   [`NOC_CONT_NOC_PORT_DATA_RANGE ]  noc__pe__port2_data            ;
  wire                                     pe__noc__port2_fc              ;
  wire   [`PE_PE_ID_BITMASK_RANGE       ]  sys__pe__port2_destinationMask ;

  // NoC port 3
  reg                                      pe__noc__port3_valid           ;
  wire   [`COMMON_STD_INTF_CNTL_RANGE ]  pe__noc__port3_cntl            ;
  wire   [`NOC_CONT_NOC_PORT_DATA_RANGE ]  pe__noc__port3_data            ;
  wire                                     noc__pe__port3_fc              ;
  wire                                     noc__pe__port3_valid           ;
  wire   [`COMMON_STD_INTF_CNTL_RANGE ]  noc__pe__port3_cntl            ;
  wire   [`NOC_CONT_NOC_PORT_DATA_RANGE ]  noc__pe__port3_data            ;
  wire                                     pe__noc__port3_fc              ;
  wire   [`PE_PE_ID_BITMASK_RANGE       ]  sys__pe__port3_destinationMask ;

