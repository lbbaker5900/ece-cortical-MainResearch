
       // Aggregate Control-Path (cp) to NoC 
      .noc__scntl__cp_ready          ( noc__scntl__cp_ready         ), 
      .scntl__noc__cp_cntl           ( scntl__noc__cp_cntl          ), 
      .scntl__noc__cp_type           ( scntl__noc__cp_type          ), 
      .scntl__noc__cp_data           ( scntl__noc__cp_data          ), 
      .scntl__noc__cp_laneId         ( scntl__noc__cp_laneId        ), 
      .scntl__noc__cp_strmId         ( scntl__noc__cp_strmId        ), 
      .scntl__noc__cp_valid          ( scntl__noc__cp_valid         ), 
       // Aggregate Data-Path (cp) from NoC 
      .scntl__noc__cp_ready          ( scntl__noc__cp_ready         ), 
      .noc__scntl__cp_cntl           ( noc__scntl__cp_cntl          ), 
      .noc__scntl__cp_type           ( noc__scntl__cp_type          ), 
      .noc__scntl__cp_data           ( noc__scntl__cp_data          ), 
      .noc__scntl__cp_peId           ( noc__scntl__cp_peId          ), 
      .noc__scntl__cp_laneId         ( noc__scntl__cp_laneId        ), 
      .noc__scntl__cp_strmId         ( noc__scntl__cp_strmId        ), 
      .noc__scntl__cp_valid          ( noc__scntl__cp_valid         ), 

       // Aggregate Data-Path (dp) to NoC 
      .noc__scntl__dp_ready          ( noc__scntl__dp_ready         ), 
      .scntl__noc__dp_cntl           ( scntl__noc__dp_cntl          ), 
      .scntl__noc__dp_type           ( scntl__noc__dp_type          ), 
      .scntl__noc__dp_peId           ( scntl__noc__dp_peId          ), 
      .scntl__noc__dp_laneId         ( scntl__noc__dp_laneId        ), 
      .scntl__noc__dp_strmId         ( scntl__noc__dp_strmId        ), 
      .scntl__noc__dp_data           ( scntl__noc__dp_data          ), 
      .scntl__noc__dp_valid          ( scntl__noc__dp_valid         ), 
       // Aggregate Data-Path (dp) from NoC 
      .scntl__noc__dp_ready          ( scntl__noc__dp_ready         ), 
      .noc__scntl__dp_cntl           ( noc__scntl__dp_cntl          ), 
      .noc__scntl__dp_type           ( noc__scntl__dp_type          ), 
      .noc__scntl__dp_laneId         ( noc__scntl__dp_laneId        ), 
      .noc__scntl__dp_strmId         ( noc__scntl__dp_strmId        ), 
      .noc__scntl__dp_data           ( noc__scntl__dp_data          ), 
      .noc__scntl__dp_valid          ( noc__scntl__dp_valid         ), 
