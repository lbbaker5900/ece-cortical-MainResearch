
            // General control and status                    
            .mgr0__sys__allSynchronized            ( mgr0__sys__allSynchronized  ),
            .sys__mgr0__thisSynchronized           ( sys__mgr0__thisSynchronized ),
            .sys__mgr0__ready                      ( sys__mgr0__ready            ),
            .sys__mgr0__complete                   ( sys__mgr0__complete         ),

            // General control and status                    
            .mgr1__sys__allSynchronized            ( mgr1__sys__allSynchronized  ),
            .sys__mgr1__thisSynchronized           ( sys__mgr1__thisSynchronized ),
            .sys__mgr1__ready                      ( sys__mgr1__ready            ),
            .sys__mgr1__complete                   ( sys__mgr1__complete         ),

            // General control and status                    
            .mgr2__sys__allSynchronized            ( mgr2__sys__allSynchronized  ),
            .sys__mgr2__thisSynchronized           ( sys__mgr2__thisSynchronized ),
            .sys__mgr2__ready                      ( sys__mgr2__ready            ),
            .sys__mgr2__complete                   ( sys__mgr2__complete         ),

            // General control and status                    
            .mgr3__sys__allSynchronized            ( mgr3__sys__allSynchronized  ),
            .sys__mgr3__thisSynchronized           ( sys__mgr3__thisSynchronized ),
            .sys__mgr3__ready                      ( sys__mgr3__ready            ),
            .sys__mgr3__complete                   ( sys__mgr3__complete         ),

            // General control and status                    
            .mgr4__sys__allSynchronized            ( mgr4__sys__allSynchronized  ),
            .sys__mgr4__thisSynchronized           ( sys__mgr4__thisSynchronized ),
            .sys__mgr4__ready                      ( sys__mgr4__ready            ),
            .sys__mgr4__complete                   ( sys__mgr4__complete         ),

            // General control and status                    
            .mgr5__sys__allSynchronized            ( mgr5__sys__allSynchronized  ),
            .sys__mgr5__thisSynchronized           ( sys__mgr5__thisSynchronized ),
            .sys__mgr5__ready                      ( sys__mgr5__ready            ),
            .sys__mgr5__complete                   ( sys__mgr5__complete         ),

            // General control and status                    
            .mgr6__sys__allSynchronized            ( mgr6__sys__allSynchronized  ),
            .sys__mgr6__thisSynchronized           ( sys__mgr6__thisSynchronized ),
            .sys__mgr6__ready                      ( sys__mgr6__ready            ),
            .sys__mgr6__complete                   ( sys__mgr6__complete         ),

            // General control and status                    
            .mgr7__sys__allSynchronized            ( mgr7__sys__allSynchronized  ),
            .sys__mgr7__thisSynchronized           ( sys__mgr7__thisSynchronized ),
            .sys__mgr7__ready                      ( sys__mgr7__ready            ),
            .sys__mgr7__complete                   ( sys__mgr7__complete         ),

            // General control and status                    
            .mgr8__sys__allSynchronized            ( mgr8__sys__allSynchronized  ),
            .sys__mgr8__thisSynchronized           ( sys__mgr8__thisSynchronized ),
            .sys__mgr8__ready                      ( sys__mgr8__ready            ),
            .sys__mgr8__complete                   ( sys__mgr8__complete         ),

            // General control and status                    
            .mgr9__sys__allSynchronized            ( mgr9__sys__allSynchronized  ),
            .sys__mgr9__thisSynchronized           ( sys__mgr9__thisSynchronized ),
            .sys__mgr9__ready                      ( sys__mgr9__ready            ),
            .sys__mgr9__complete                   ( sys__mgr9__complete         ),

            // General control and status                    
            .mgr10__sys__allSynchronized            ( mgr10__sys__allSynchronized  ),
            .sys__mgr10__thisSynchronized           ( sys__mgr10__thisSynchronized ),
            .sys__mgr10__ready                      ( sys__mgr10__ready            ),
            .sys__mgr10__complete                   ( sys__mgr10__complete         ),

            // General control and status                    
            .mgr11__sys__allSynchronized            ( mgr11__sys__allSynchronized  ),
            .sys__mgr11__thisSynchronized           ( sys__mgr11__thisSynchronized ),
            .sys__mgr11__ready                      ( sys__mgr11__ready            ),
            .sys__mgr11__complete                   ( sys__mgr11__complete         ),

            // General control and status                    
            .mgr12__sys__allSynchronized            ( mgr12__sys__allSynchronized  ),
            .sys__mgr12__thisSynchronized           ( sys__mgr12__thisSynchronized ),
            .sys__mgr12__ready                      ( sys__mgr12__ready            ),
            .sys__mgr12__complete                   ( sys__mgr12__complete         ),

            // General control and status                    
            .mgr13__sys__allSynchronized            ( mgr13__sys__allSynchronized  ),
            .sys__mgr13__thisSynchronized           ( sys__mgr13__thisSynchronized ),
            .sys__mgr13__ready                      ( sys__mgr13__ready            ),
            .sys__mgr13__complete                   ( sys__mgr13__complete         ),

            // General control and status                    
            .mgr14__sys__allSynchronized            ( mgr14__sys__allSynchronized  ),
            .sys__mgr14__thisSynchronized           ( sys__mgr14__thisSynchronized ),
            .sys__mgr14__ready                      ( sys__mgr14__ready            ),
            .sys__mgr14__complete                   ( sys__mgr14__complete         ),

            // General control and status                    
            .mgr15__sys__allSynchronized            ( mgr15__sys__allSynchronized  ),
            .sys__mgr15__thisSynchronized           ( sys__mgr15__thisSynchronized ),
            .sys__mgr15__ready                      ( sys__mgr15__ready            ),
            .sys__mgr15__complete                   ( sys__mgr15__complete         ),

            // General control and status                    
            .mgr16__sys__allSynchronized            ( mgr16__sys__allSynchronized  ),
            .sys__mgr16__thisSynchronized           ( sys__mgr16__thisSynchronized ),
            .sys__mgr16__ready                      ( sys__mgr16__ready            ),
            .sys__mgr16__complete                   ( sys__mgr16__complete         ),

            // General control and status                    
            .mgr17__sys__allSynchronized            ( mgr17__sys__allSynchronized  ),
            .sys__mgr17__thisSynchronized           ( sys__mgr17__thisSynchronized ),
            .sys__mgr17__ready                      ( sys__mgr17__ready            ),
            .sys__mgr17__complete                   ( sys__mgr17__complete         ),

            // General control and status                    
            .mgr18__sys__allSynchronized            ( mgr18__sys__allSynchronized  ),
            .sys__mgr18__thisSynchronized           ( sys__mgr18__thisSynchronized ),
            .sys__mgr18__ready                      ( sys__mgr18__ready            ),
            .sys__mgr18__complete                   ( sys__mgr18__complete         ),

            // General control and status                    
            .mgr19__sys__allSynchronized            ( mgr19__sys__allSynchronized  ),
            .sys__mgr19__thisSynchronized           ( sys__mgr19__thisSynchronized ),
            .sys__mgr19__ready                      ( sys__mgr19__ready            ),
            .sys__mgr19__complete                   ( sys__mgr19__complete         ),

            // General control and status                    
            .mgr20__sys__allSynchronized            ( mgr20__sys__allSynchronized  ),
            .sys__mgr20__thisSynchronized           ( sys__mgr20__thisSynchronized ),
            .sys__mgr20__ready                      ( sys__mgr20__ready            ),
            .sys__mgr20__complete                   ( sys__mgr20__complete         ),

            // General control and status                    
            .mgr21__sys__allSynchronized            ( mgr21__sys__allSynchronized  ),
            .sys__mgr21__thisSynchronized           ( sys__mgr21__thisSynchronized ),
            .sys__mgr21__ready                      ( sys__mgr21__ready            ),
            .sys__mgr21__complete                   ( sys__mgr21__complete         ),

            // General control and status                    
            .mgr22__sys__allSynchronized            ( mgr22__sys__allSynchronized  ),
            .sys__mgr22__thisSynchronized           ( sys__mgr22__thisSynchronized ),
            .sys__mgr22__ready                      ( sys__mgr22__ready            ),
            .sys__mgr22__complete                   ( sys__mgr22__complete         ),

            // General control and status                    
            .mgr23__sys__allSynchronized            ( mgr23__sys__allSynchronized  ),
            .sys__mgr23__thisSynchronized           ( sys__mgr23__thisSynchronized ),
            .sys__mgr23__ready                      ( sys__mgr23__ready            ),
            .sys__mgr23__complete                   ( sys__mgr23__complete         ),

            // General control and status                    
            .mgr24__sys__allSynchronized            ( mgr24__sys__allSynchronized  ),
            .sys__mgr24__thisSynchronized           ( sys__mgr24__thisSynchronized ),
            .sys__mgr24__ready                      ( sys__mgr24__ready            ),
            .sys__mgr24__complete                   ( sys__mgr24__complete         ),

            // General control and status                    
            .mgr25__sys__allSynchronized            ( mgr25__sys__allSynchronized  ),
            .sys__mgr25__thisSynchronized           ( sys__mgr25__thisSynchronized ),
            .sys__mgr25__ready                      ( sys__mgr25__ready            ),
            .sys__mgr25__complete                   ( sys__mgr25__complete         ),

            // General control and status                    
            .mgr26__sys__allSynchronized            ( mgr26__sys__allSynchronized  ),
            .sys__mgr26__thisSynchronized           ( sys__mgr26__thisSynchronized ),
            .sys__mgr26__ready                      ( sys__mgr26__ready            ),
            .sys__mgr26__complete                   ( sys__mgr26__complete         ),

            // General control and status                    
            .mgr27__sys__allSynchronized            ( mgr27__sys__allSynchronized  ),
            .sys__mgr27__thisSynchronized           ( sys__mgr27__thisSynchronized ),
            .sys__mgr27__ready                      ( sys__mgr27__ready            ),
            .sys__mgr27__complete                   ( sys__mgr27__complete         ),

            // General control and status                    
            .mgr28__sys__allSynchronized            ( mgr28__sys__allSynchronized  ),
            .sys__mgr28__thisSynchronized           ( sys__mgr28__thisSynchronized ),
            .sys__mgr28__ready                      ( sys__mgr28__ready            ),
            .sys__mgr28__complete                   ( sys__mgr28__complete         ),

            // General control and status                    
            .mgr29__sys__allSynchronized            ( mgr29__sys__allSynchronized  ),
            .sys__mgr29__thisSynchronized           ( sys__mgr29__thisSynchronized ),
            .sys__mgr29__ready                      ( sys__mgr29__ready            ),
            .sys__mgr29__complete                   ( sys__mgr29__complete         ),

            // General control and status                    
            .mgr30__sys__allSynchronized            ( mgr30__sys__allSynchronized  ),
            .sys__mgr30__thisSynchronized           ( sys__mgr30__thisSynchronized ),
            .sys__mgr30__ready                      ( sys__mgr30__ready            ),
            .sys__mgr30__complete                   ( sys__mgr30__complete         ),

            // General control and status                    
            .mgr31__sys__allSynchronized            ( mgr31__sys__allSynchronized  ),
            .sys__mgr31__thisSynchronized           ( sys__mgr31__thisSynchronized ),
            .sys__mgr31__ready                      ( sys__mgr31__ready            ),
            .sys__mgr31__complete                   ( sys__mgr31__complete         ),

            // General control and status                    
            .mgr32__sys__allSynchronized            ( mgr32__sys__allSynchronized  ),
            .sys__mgr32__thisSynchronized           ( sys__mgr32__thisSynchronized ),
            .sys__mgr32__ready                      ( sys__mgr32__ready            ),
            .sys__mgr32__complete                   ( sys__mgr32__complete         ),

            // General control and status                    
            .mgr33__sys__allSynchronized            ( mgr33__sys__allSynchronized  ),
            .sys__mgr33__thisSynchronized           ( sys__mgr33__thisSynchronized ),
            .sys__mgr33__ready                      ( sys__mgr33__ready            ),
            .sys__mgr33__complete                   ( sys__mgr33__complete         ),

            // General control and status                    
            .mgr34__sys__allSynchronized            ( mgr34__sys__allSynchronized  ),
            .sys__mgr34__thisSynchronized           ( sys__mgr34__thisSynchronized ),
            .sys__mgr34__ready                      ( sys__mgr34__ready            ),
            .sys__mgr34__complete                   ( sys__mgr34__complete         ),

            // General control and status                    
            .mgr35__sys__allSynchronized            ( mgr35__sys__allSynchronized  ),
            .sys__mgr35__thisSynchronized           ( sys__mgr35__thisSynchronized ),
            .sys__mgr35__ready                      ( sys__mgr35__ready            ),
            .sys__mgr35__complete                   ( sys__mgr35__complete         ),

            // General control and status                    
            .mgr36__sys__allSynchronized            ( mgr36__sys__allSynchronized  ),
            .sys__mgr36__thisSynchronized           ( sys__mgr36__thisSynchronized ),
            .sys__mgr36__ready                      ( sys__mgr36__ready            ),
            .sys__mgr36__complete                   ( sys__mgr36__complete         ),

            // General control and status                    
            .mgr37__sys__allSynchronized            ( mgr37__sys__allSynchronized  ),
            .sys__mgr37__thisSynchronized           ( sys__mgr37__thisSynchronized ),
            .sys__mgr37__ready                      ( sys__mgr37__ready            ),
            .sys__mgr37__complete                   ( sys__mgr37__complete         ),

            // General control and status                    
            .mgr38__sys__allSynchronized            ( mgr38__sys__allSynchronized  ),
            .sys__mgr38__thisSynchronized           ( sys__mgr38__thisSynchronized ),
            .sys__mgr38__ready                      ( sys__mgr38__ready            ),
            .sys__mgr38__complete                   ( sys__mgr38__complete         ),

            // General control and status                    
            .mgr39__sys__allSynchronized            ( mgr39__sys__allSynchronized  ),
            .sys__mgr39__thisSynchronized           ( sys__mgr39__thisSynchronized ),
            .sys__mgr39__ready                      ( sys__mgr39__ready            ),
            .sys__mgr39__complete                   ( sys__mgr39__complete         ),

            // General control and status                    
            .mgr40__sys__allSynchronized            ( mgr40__sys__allSynchronized  ),
            .sys__mgr40__thisSynchronized           ( sys__mgr40__thisSynchronized ),
            .sys__mgr40__ready                      ( sys__mgr40__ready            ),
            .sys__mgr40__complete                   ( sys__mgr40__complete         ),

            // General control and status                    
            .mgr41__sys__allSynchronized            ( mgr41__sys__allSynchronized  ),
            .sys__mgr41__thisSynchronized           ( sys__mgr41__thisSynchronized ),
            .sys__mgr41__ready                      ( sys__mgr41__ready            ),
            .sys__mgr41__complete                   ( sys__mgr41__complete         ),

            // General control and status                    
            .mgr42__sys__allSynchronized            ( mgr42__sys__allSynchronized  ),
            .sys__mgr42__thisSynchronized           ( sys__mgr42__thisSynchronized ),
            .sys__mgr42__ready                      ( sys__mgr42__ready            ),
            .sys__mgr42__complete                   ( sys__mgr42__complete         ),

            // General control and status                    
            .mgr43__sys__allSynchronized            ( mgr43__sys__allSynchronized  ),
            .sys__mgr43__thisSynchronized           ( sys__mgr43__thisSynchronized ),
            .sys__mgr43__ready                      ( sys__mgr43__ready            ),
            .sys__mgr43__complete                   ( sys__mgr43__complete         ),

            // General control and status                    
            .mgr44__sys__allSynchronized            ( mgr44__sys__allSynchronized  ),
            .sys__mgr44__thisSynchronized           ( sys__mgr44__thisSynchronized ),
            .sys__mgr44__ready                      ( sys__mgr44__ready            ),
            .sys__mgr44__complete                   ( sys__mgr44__complete         ),

            // General control and status                    
            .mgr45__sys__allSynchronized            ( mgr45__sys__allSynchronized  ),
            .sys__mgr45__thisSynchronized           ( sys__mgr45__thisSynchronized ),
            .sys__mgr45__ready                      ( sys__mgr45__ready            ),
            .sys__mgr45__complete                   ( sys__mgr45__complete         ),

            // General control and status                    
            .mgr46__sys__allSynchronized            ( mgr46__sys__allSynchronized  ),
            .sys__mgr46__thisSynchronized           ( sys__mgr46__thisSynchronized ),
            .sys__mgr46__ready                      ( sys__mgr46__ready            ),
            .sys__mgr46__complete                   ( sys__mgr46__complete         ),

            // General control and status                    
            .mgr47__sys__allSynchronized            ( mgr47__sys__allSynchronized  ),
            .sys__mgr47__thisSynchronized           ( sys__mgr47__thisSynchronized ),
            .sys__mgr47__ready                      ( sys__mgr47__ready            ),
            .sys__mgr47__complete                   ( sys__mgr47__complete         ),

            // General control and status                    
            .mgr48__sys__allSynchronized            ( mgr48__sys__allSynchronized  ),
            .sys__mgr48__thisSynchronized           ( sys__mgr48__thisSynchronized ),
            .sys__mgr48__ready                      ( sys__mgr48__ready            ),
            .sys__mgr48__complete                   ( sys__mgr48__complete         ),

            // General control and status                    
            .mgr49__sys__allSynchronized            ( mgr49__sys__allSynchronized  ),
            .sys__mgr49__thisSynchronized           ( sys__mgr49__thisSynchronized ),
            .sys__mgr49__ready                      ( sys__mgr49__ready            ),
            .sys__mgr49__complete                   ( sys__mgr49__complete         ),

            // General control and status                    
            .mgr50__sys__allSynchronized            ( mgr50__sys__allSynchronized  ),
            .sys__mgr50__thisSynchronized           ( sys__mgr50__thisSynchronized ),
            .sys__mgr50__ready                      ( sys__mgr50__ready            ),
            .sys__mgr50__complete                   ( sys__mgr50__complete         ),

            // General control and status                    
            .mgr51__sys__allSynchronized            ( mgr51__sys__allSynchronized  ),
            .sys__mgr51__thisSynchronized           ( sys__mgr51__thisSynchronized ),
            .sys__mgr51__ready                      ( sys__mgr51__ready            ),
            .sys__mgr51__complete                   ( sys__mgr51__complete         ),

            // General control and status                    
            .mgr52__sys__allSynchronized            ( mgr52__sys__allSynchronized  ),
            .sys__mgr52__thisSynchronized           ( sys__mgr52__thisSynchronized ),
            .sys__mgr52__ready                      ( sys__mgr52__ready            ),
            .sys__mgr52__complete                   ( sys__mgr52__complete         ),

            // General control and status                    
            .mgr53__sys__allSynchronized            ( mgr53__sys__allSynchronized  ),
            .sys__mgr53__thisSynchronized           ( sys__mgr53__thisSynchronized ),
            .sys__mgr53__ready                      ( sys__mgr53__ready            ),
            .sys__mgr53__complete                   ( sys__mgr53__complete         ),

            // General control and status                    
            .mgr54__sys__allSynchronized            ( mgr54__sys__allSynchronized  ),
            .sys__mgr54__thisSynchronized           ( sys__mgr54__thisSynchronized ),
            .sys__mgr54__ready                      ( sys__mgr54__ready            ),
            .sys__mgr54__complete                   ( sys__mgr54__complete         ),

            // General control and status                    
            .mgr55__sys__allSynchronized            ( mgr55__sys__allSynchronized  ),
            .sys__mgr55__thisSynchronized           ( sys__mgr55__thisSynchronized ),
            .sys__mgr55__ready                      ( sys__mgr55__ready            ),
            .sys__mgr55__complete                   ( sys__mgr55__complete         ),

            // General control and status                    
            .mgr56__sys__allSynchronized            ( mgr56__sys__allSynchronized  ),
            .sys__mgr56__thisSynchronized           ( sys__mgr56__thisSynchronized ),
            .sys__mgr56__ready                      ( sys__mgr56__ready            ),
            .sys__mgr56__complete                   ( sys__mgr56__complete         ),

            // General control and status                    
            .mgr57__sys__allSynchronized            ( mgr57__sys__allSynchronized  ),
            .sys__mgr57__thisSynchronized           ( sys__mgr57__thisSynchronized ),
            .sys__mgr57__ready                      ( sys__mgr57__ready            ),
            .sys__mgr57__complete                   ( sys__mgr57__complete         ),

            // General control and status                    
            .mgr58__sys__allSynchronized            ( mgr58__sys__allSynchronized  ),
            .sys__mgr58__thisSynchronized           ( sys__mgr58__thisSynchronized ),
            .sys__mgr58__ready                      ( sys__mgr58__ready            ),
            .sys__mgr58__complete                   ( sys__mgr58__complete         ),

            // General control and status                    
            .mgr59__sys__allSynchronized            ( mgr59__sys__allSynchronized  ),
            .sys__mgr59__thisSynchronized           ( sys__mgr59__thisSynchronized ),
            .sys__mgr59__ready                      ( sys__mgr59__ready            ),
            .sys__mgr59__complete                   ( sys__mgr59__complete         ),

            // General control and status                    
            .mgr60__sys__allSynchronized            ( mgr60__sys__allSynchronized  ),
            .sys__mgr60__thisSynchronized           ( sys__mgr60__thisSynchronized ),
            .sys__mgr60__ready                      ( sys__mgr60__ready            ),
            .sys__mgr60__complete                   ( sys__mgr60__complete         ),

            // General control and status                    
            .mgr61__sys__allSynchronized            ( mgr61__sys__allSynchronized  ),
            .sys__mgr61__thisSynchronized           ( sys__mgr61__thisSynchronized ),
            .sys__mgr61__ready                      ( sys__mgr61__ready            ),
            .sys__mgr61__complete                   ( sys__mgr61__complete         ),

            // General control and status                    
            .mgr62__sys__allSynchronized            ( mgr62__sys__allSynchronized  ),
            .sys__mgr62__thisSynchronized           ( sys__mgr62__thisSynchronized ),
            .sys__mgr62__ready                      ( sys__mgr62__ready            ),
            .sys__mgr62__complete                   ( sys__mgr62__complete         ),

            // General control and status                    
            .mgr63__sys__allSynchronized            ( mgr63__sys__allSynchronized  ),
            .sys__mgr63__thisSynchronized           ( sys__mgr63__thisSynchronized ),
            .sys__mgr63__ready                      ( sys__mgr63__ready            ),
            .sys__mgr63__complete                   ( sys__mgr63__complete         ),
