
               // Lane 0                 
               .pe__std__lane0_strm0_ready         ( pe__std__lane0_strm0_ready      ),      
               .std__pe__lane0_strm0_cntl          ( std__pe__lane0_strm0_cntl       ),      
               .std__pe__lane0_strm0_data          ( std__pe__lane0_strm0_data       ),      
               .std__pe__lane0_strm0_data_valid    ( std__pe__lane0_strm0_data_valid ),      
               .std__pe__lane0_strm0_data_mask     ( std__pe__lane0_strm0_data_mask  ),      
               .pe__std__lane0_strm1_ready         ( pe__std__lane0_strm1_ready      ),      
               .std__pe__lane0_strm1_cntl          ( std__pe__lane0_strm1_cntl       ),      
               .std__pe__lane0_strm1_data          ( std__pe__lane0_strm1_data       ),      
               .std__pe__lane0_strm1_data_valid    ( std__pe__lane0_strm1_data_valid ),      
               .std__pe__lane0_strm1_data_mask     ( std__pe__lane0_strm1_data_mask  ),      
               // Lane 1                 
               .pe__std__lane1_strm0_ready         ( pe__std__lane1_strm0_ready      ),      
               .std__pe__lane1_strm0_cntl          ( std__pe__lane1_strm0_cntl       ),      
               .std__pe__lane1_strm0_data          ( std__pe__lane1_strm0_data       ),      
               .std__pe__lane1_strm0_data_valid    ( std__pe__lane1_strm0_data_valid ),      
               .std__pe__lane1_strm0_data_mask     ( std__pe__lane1_strm0_data_mask  ),      
               .pe__std__lane1_strm1_ready         ( pe__std__lane1_strm1_ready      ),      
               .std__pe__lane1_strm1_cntl          ( std__pe__lane1_strm1_cntl       ),      
               .std__pe__lane1_strm1_data          ( std__pe__lane1_strm1_data       ),      
               .std__pe__lane1_strm1_data_valid    ( std__pe__lane1_strm1_data_valid ),      
               .std__pe__lane1_strm1_data_mask     ( std__pe__lane1_strm1_data_mask  ),      
               // Lane 2                 
               .pe__std__lane2_strm0_ready         ( pe__std__lane2_strm0_ready      ),      
               .std__pe__lane2_strm0_cntl          ( std__pe__lane2_strm0_cntl       ),      
               .std__pe__lane2_strm0_data          ( std__pe__lane2_strm0_data       ),      
               .std__pe__lane2_strm0_data_valid    ( std__pe__lane2_strm0_data_valid ),      
               .std__pe__lane2_strm0_data_mask     ( std__pe__lane2_strm0_data_mask  ),      
               .pe__std__lane2_strm1_ready         ( pe__std__lane2_strm1_ready      ),      
               .std__pe__lane2_strm1_cntl          ( std__pe__lane2_strm1_cntl       ),      
               .std__pe__lane2_strm1_data          ( std__pe__lane2_strm1_data       ),      
               .std__pe__lane2_strm1_data_valid    ( std__pe__lane2_strm1_data_valid ),      
               .std__pe__lane2_strm1_data_mask     ( std__pe__lane2_strm1_data_mask  ),      
               // Lane 3                 
               .pe__std__lane3_strm0_ready         ( pe__std__lane3_strm0_ready      ),      
               .std__pe__lane3_strm0_cntl          ( std__pe__lane3_strm0_cntl       ),      
               .std__pe__lane3_strm0_data          ( std__pe__lane3_strm0_data       ),      
               .std__pe__lane3_strm0_data_valid    ( std__pe__lane3_strm0_data_valid ),      
               .std__pe__lane3_strm0_data_mask     ( std__pe__lane3_strm0_data_mask  ),      
               .pe__std__lane3_strm1_ready         ( pe__std__lane3_strm1_ready      ),      
               .std__pe__lane3_strm1_cntl          ( std__pe__lane3_strm1_cntl       ),      
               .std__pe__lane3_strm1_data          ( std__pe__lane3_strm1_data       ),      
               .std__pe__lane3_strm1_data_valid    ( std__pe__lane3_strm1_data_valid ),      
               .std__pe__lane3_strm1_data_mask     ( std__pe__lane3_strm1_data_mask  ),      
               // Lane 4                 
               .pe__std__lane4_strm0_ready         ( pe__std__lane4_strm0_ready      ),      
               .std__pe__lane4_strm0_cntl          ( std__pe__lane4_strm0_cntl       ),      
               .std__pe__lane4_strm0_data          ( std__pe__lane4_strm0_data       ),      
               .std__pe__lane4_strm0_data_valid    ( std__pe__lane4_strm0_data_valid ),      
               .std__pe__lane4_strm0_data_mask     ( std__pe__lane4_strm0_data_mask  ),      
               .pe__std__lane4_strm1_ready         ( pe__std__lane4_strm1_ready      ),      
               .std__pe__lane4_strm1_cntl          ( std__pe__lane4_strm1_cntl       ),      
               .std__pe__lane4_strm1_data          ( std__pe__lane4_strm1_data       ),      
               .std__pe__lane4_strm1_data_valid    ( std__pe__lane4_strm1_data_valid ),      
               .std__pe__lane4_strm1_data_mask     ( std__pe__lane4_strm1_data_mask  ),      
               // Lane 5                 
               .pe__std__lane5_strm0_ready         ( pe__std__lane5_strm0_ready      ),      
               .std__pe__lane5_strm0_cntl          ( std__pe__lane5_strm0_cntl       ),      
               .std__pe__lane5_strm0_data          ( std__pe__lane5_strm0_data       ),      
               .std__pe__lane5_strm0_data_valid    ( std__pe__lane5_strm0_data_valid ),      
               .std__pe__lane5_strm0_data_mask     ( std__pe__lane5_strm0_data_mask  ),      
               .pe__std__lane5_strm1_ready         ( pe__std__lane5_strm1_ready      ),      
               .std__pe__lane5_strm1_cntl          ( std__pe__lane5_strm1_cntl       ),      
               .std__pe__lane5_strm1_data          ( std__pe__lane5_strm1_data       ),      
               .std__pe__lane5_strm1_data_valid    ( std__pe__lane5_strm1_data_valid ),      
               .std__pe__lane5_strm1_data_mask     ( std__pe__lane5_strm1_data_mask  ),      
               // Lane 6                 
               .pe__std__lane6_strm0_ready         ( pe__std__lane6_strm0_ready      ),      
               .std__pe__lane6_strm0_cntl          ( std__pe__lane6_strm0_cntl       ),      
               .std__pe__lane6_strm0_data          ( std__pe__lane6_strm0_data       ),      
               .std__pe__lane6_strm0_data_valid    ( std__pe__lane6_strm0_data_valid ),      
               .std__pe__lane6_strm0_data_mask     ( std__pe__lane6_strm0_data_mask  ),      
               .pe__std__lane6_strm1_ready         ( pe__std__lane6_strm1_ready      ),      
               .std__pe__lane6_strm1_cntl          ( std__pe__lane6_strm1_cntl       ),      
               .std__pe__lane6_strm1_data          ( std__pe__lane6_strm1_data       ),      
               .std__pe__lane6_strm1_data_valid    ( std__pe__lane6_strm1_data_valid ),      
               .std__pe__lane6_strm1_data_mask     ( std__pe__lane6_strm1_data_mask  ),      
               // Lane 7                 
               .pe__std__lane7_strm0_ready         ( pe__std__lane7_strm0_ready      ),      
               .std__pe__lane7_strm0_cntl          ( std__pe__lane7_strm0_cntl       ),      
               .std__pe__lane7_strm0_data          ( std__pe__lane7_strm0_data       ),      
               .std__pe__lane7_strm0_data_valid    ( std__pe__lane7_strm0_data_valid ),      
               .std__pe__lane7_strm0_data_mask     ( std__pe__lane7_strm0_data_mask  ),      
               .pe__std__lane7_strm1_ready         ( pe__std__lane7_strm1_ready      ),      
               .std__pe__lane7_strm1_cntl          ( std__pe__lane7_strm1_cntl       ),      
               .std__pe__lane7_strm1_data          ( std__pe__lane7_strm1_data       ),      
               .std__pe__lane7_strm1_data_valid    ( std__pe__lane7_strm1_data_valid ),      
               .std__pe__lane7_strm1_data_mask     ( std__pe__lane7_strm1_data_mask  ),      
               // Lane 8                 
               .pe__std__lane8_strm0_ready         ( pe__std__lane8_strm0_ready      ),      
               .std__pe__lane8_strm0_cntl          ( std__pe__lane8_strm0_cntl       ),      
               .std__pe__lane8_strm0_data          ( std__pe__lane8_strm0_data       ),      
               .std__pe__lane8_strm0_data_valid    ( std__pe__lane8_strm0_data_valid ),      
               .std__pe__lane8_strm0_data_mask     ( std__pe__lane8_strm0_data_mask  ),      
               .pe__std__lane8_strm1_ready         ( pe__std__lane8_strm1_ready      ),      
               .std__pe__lane8_strm1_cntl          ( std__pe__lane8_strm1_cntl       ),      
               .std__pe__lane8_strm1_data          ( std__pe__lane8_strm1_data       ),      
               .std__pe__lane8_strm1_data_valid    ( std__pe__lane8_strm1_data_valid ),      
               .std__pe__lane8_strm1_data_mask     ( std__pe__lane8_strm1_data_mask  ),      
               // Lane 9                 
               .pe__std__lane9_strm0_ready         ( pe__std__lane9_strm0_ready      ),      
               .std__pe__lane9_strm0_cntl          ( std__pe__lane9_strm0_cntl       ),      
               .std__pe__lane9_strm0_data          ( std__pe__lane9_strm0_data       ),      
               .std__pe__lane9_strm0_data_valid    ( std__pe__lane9_strm0_data_valid ),      
               .std__pe__lane9_strm0_data_mask     ( std__pe__lane9_strm0_data_mask  ),      
               .pe__std__lane9_strm1_ready         ( pe__std__lane9_strm1_ready      ),      
               .std__pe__lane9_strm1_cntl          ( std__pe__lane9_strm1_cntl       ),      
               .std__pe__lane9_strm1_data          ( std__pe__lane9_strm1_data       ),      
               .std__pe__lane9_strm1_data_valid    ( std__pe__lane9_strm1_data_valid ),      
               .std__pe__lane9_strm1_data_mask     ( std__pe__lane9_strm1_data_mask  ),      
               // Lane 10                 
               .pe__std__lane10_strm0_ready         ( pe__std__lane10_strm0_ready      ),      
               .std__pe__lane10_strm0_cntl          ( std__pe__lane10_strm0_cntl       ),      
               .std__pe__lane10_strm0_data          ( std__pe__lane10_strm0_data       ),      
               .std__pe__lane10_strm0_data_valid    ( std__pe__lane10_strm0_data_valid ),      
               .std__pe__lane10_strm0_data_mask     ( std__pe__lane10_strm0_data_mask  ),      
               .pe__std__lane10_strm1_ready         ( pe__std__lane10_strm1_ready      ),      
               .std__pe__lane10_strm1_cntl          ( std__pe__lane10_strm1_cntl       ),      
               .std__pe__lane10_strm1_data          ( std__pe__lane10_strm1_data       ),      
               .std__pe__lane10_strm1_data_valid    ( std__pe__lane10_strm1_data_valid ),      
               .std__pe__lane10_strm1_data_mask     ( std__pe__lane10_strm1_data_mask  ),      
               // Lane 11                 
               .pe__std__lane11_strm0_ready         ( pe__std__lane11_strm0_ready      ),      
               .std__pe__lane11_strm0_cntl          ( std__pe__lane11_strm0_cntl       ),      
               .std__pe__lane11_strm0_data          ( std__pe__lane11_strm0_data       ),      
               .std__pe__lane11_strm0_data_valid    ( std__pe__lane11_strm0_data_valid ),      
               .std__pe__lane11_strm0_data_mask     ( std__pe__lane11_strm0_data_mask  ),      
               .pe__std__lane11_strm1_ready         ( pe__std__lane11_strm1_ready      ),      
               .std__pe__lane11_strm1_cntl          ( std__pe__lane11_strm1_cntl       ),      
               .std__pe__lane11_strm1_data          ( std__pe__lane11_strm1_data       ),      
               .std__pe__lane11_strm1_data_valid    ( std__pe__lane11_strm1_data_valid ),      
               .std__pe__lane11_strm1_data_mask     ( std__pe__lane11_strm1_data_mask  ),      
               // Lane 12                 
               .pe__std__lane12_strm0_ready         ( pe__std__lane12_strm0_ready      ),      
               .std__pe__lane12_strm0_cntl          ( std__pe__lane12_strm0_cntl       ),      
               .std__pe__lane12_strm0_data          ( std__pe__lane12_strm0_data       ),      
               .std__pe__lane12_strm0_data_valid    ( std__pe__lane12_strm0_data_valid ),      
               .std__pe__lane12_strm0_data_mask     ( std__pe__lane12_strm0_data_mask  ),      
               .pe__std__lane12_strm1_ready         ( pe__std__lane12_strm1_ready      ),      
               .std__pe__lane12_strm1_cntl          ( std__pe__lane12_strm1_cntl       ),      
               .std__pe__lane12_strm1_data          ( std__pe__lane12_strm1_data       ),      
               .std__pe__lane12_strm1_data_valid    ( std__pe__lane12_strm1_data_valid ),      
               .std__pe__lane12_strm1_data_mask     ( std__pe__lane12_strm1_data_mask  ),      
               // Lane 13                 
               .pe__std__lane13_strm0_ready         ( pe__std__lane13_strm0_ready      ),      
               .std__pe__lane13_strm0_cntl          ( std__pe__lane13_strm0_cntl       ),      
               .std__pe__lane13_strm0_data          ( std__pe__lane13_strm0_data       ),      
               .std__pe__lane13_strm0_data_valid    ( std__pe__lane13_strm0_data_valid ),      
               .std__pe__lane13_strm0_data_mask     ( std__pe__lane13_strm0_data_mask  ),      
               .pe__std__lane13_strm1_ready         ( pe__std__lane13_strm1_ready      ),      
               .std__pe__lane13_strm1_cntl          ( std__pe__lane13_strm1_cntl       ),      
               .std__pe__lane13_strm1_data          ( std__pe__lane13_strm1_data       ),      
               .std__pe__lane13_strm1_data_valid    ( std__pe__lane13_strm1_data_valid ),      
               .std__pe__lane13_strm1_data_mask     ( std__pe__lane13_strm1_data_mask  ),      
               // Lane 14                 
               .pe__std__lane14_strm0_ready         ( pe__std__lane14_strm0_ready      ),      
               .std__pe__lane14_strm0_cntl          ( std__pe__lane14_strm0_cntl       ),      
               .std__pe__lane14_strm0_data          ( std__pe__lane14_strm0_data       ),      
               .std__pe__lane14_strm0_data_valid    ( std__pe__lane14_strm0_data_valid ),      
               .std__pe__lane14_strm0_data_mask     ( std__pe__lane14_strm0_data_mask  ),      
               .pe__std__lane14_strm1_ready         ( pe__std__lane14_strm1_ready      ),      
               .std__pe__lane14_strm1_cntl          ( std__pe__lane14_strm1_cntl       ),      
               .std__pe__lane14_strm1_data          ( std__pe__lane14_strm1_data       ),      
               .std__pe__lane14_strm1_data_valid    ( std__pe__lane14_strm1_data_valid ),      
               .std__pe__lane14_strm1_data_mask     ( std__pe__lane14_strm1_data_mask  ),      
               // Lane 15                 
               .pe__std__lane15_strm0_ready         ( pe__std__lane15_strm0_ready      ),      
               .std__pe__lane15_strm0_cntl          ( std__pe__lane15_strm0_cntl       ),      
               .std__pe__lane15_strm0_data          ( std__pe__lane15_strm0_data       ),      
               .std__pe__lane15_strm0_data_valid    ( std__pe__lane15_strm0_data_valid ),      
               .std__pe__lane15_strm0_data_mask     ( std__pe__lane15_strm0_data_mask  ),      
               .pe__std__lane15_strm1_ready         ( pe__std__lane15_strm1_ready      ),      
               .std__pe__lane15_strm1_cntl          ( std__pe__lane15_strm1_cntl       ),      
               .std__pe__lane15_strm1_data          ( std__pe__lane15_strm1_data       ),      
               .std__pe__lane15_strm1_data_valid    ( std__pe__lane15_strm1_data_valid ),      
               .std__pe__lane15_strm1_data_mask     ( std__pe__lane15_strm1_data_mask  ),      
               // Lane 16                 
               .pe__std__lane16_strm0_ready         ( pe__std__lane16_strm0_ready      ),      
               .std__pe__lane16_strm0_cntl          ( std__pe__lane16_strm0_cntl       ),      
               .std__pe__lane16_strm0_data          ( std__pe__lane16_strm0_data       ),      
               .std__pe__lane16_strm0_data_valid    ( std__pe__lane16_strm0_data_valid ),      
               .std__pe__lane16_strm0_data_mask     ( std__pe__lane16_strm0_data_mask  ),      
               .pe__std__lane16_strm1_ready         ( pe__std__lane16_strm1_ready      ),      
               .std__pe__lane16_strm1_cntl          ( std__pe__lane16_strm1_cntl       ),      
               .std__pe__lane16_strm1_data          ( std__pe__lane16_strm1_data       ),      
               .std__pe__lane16_strm1_data_valid    ( std__pe__lane16_strm1_data_valid ),      
               .std__pe__lane16_strm1_data_mask     ( std__pe__lane16_strm1_data_mask  ),      
               // Lane 17                 
               .pe__std__lane17_strm0_ready         ( pe__std__lane17_strm0_ready      ),      
               .std__pe__lane17_strm0_cntl          ( std__pe__lane17_strm0_cntl       ),      
               .std__pe__lane17_strm0_data          ( std__pe__lane17_strm0_data       ),      
               .std__pe__lane17_strm0_data_valid    ( std__pe__lane17_strm0_data_valid ),      
               .std__pe__lane17_strm0_data_mask     ( std__pe__lane17_strm0_data_mask  ),      
               .pe__std__lane17_strm1_ready         ( pe__std__lane17_strm1_ready      ),      
               .std__pe__lane17_strm1_cntl          ( std__pe__lane17_strm1_cntl       ),      
               .std__pe__lane17_strm1_data          ( std__pe__lane17_strm1_data       ),      
               .std__pe__lane17_strm1_data_valid    ( std__pe__lane17_strm1_data_valid ),      
               .std__pe__lane17_strm1_data_mask     ( std__pe__lane17_strm1_data_mask  ),      
               // Lane 18                 
               .pe__std__lane18_strm0_ready         ( pe__std__lane18_strm0_ready      ),      
               .std__pe__lane18_strm0_cntl          ( std__pe__lane18_strm0_cntl       ),      
               .std__pe__lane18_strm0_data          ( std__pe__lane18_strm0_data       ),      
               .std__pe__lane18_strm0_data_valid    ( std__pe__lane18_strm0_data_valid ),      
               .std__pe__lane18_strm0_data_mask     ( std__pe__lane18_strm0_data_mask  ),      
               .pe__std__lane18_strm1_ready         ( pe__std__lane18_strm1_ready      ),      
               .std__pe__lane18_strm1_cntl          ( std__pe__lane18_strm1_cntl       ),      
               .std__pe__lane18_strm1_data          ( std__pe__lane18_strm1_data       ),      
               .std__pe__lane18_strm1_data_valid    ( std__pe__lane18_strm1_data_valid ),      
               .std__pe__lane18_strm1_data_mask     ( std__pe__lane18_strm1_data_mask  ),      
               // Lane 19                 
               .pe__std__lane19_strm0_ready         ( pe__std__lane19_strm0_ready      ),      
               .std__pe__lane19_strm0_cntl          ( std__pe__lane19_strm0_cntl       ),      
               .std__pe__lane19_strm0_data          ( std__pe__lane19_strm0_data       ),      
               .std__pe__lane19_strm0_data_valid    ( std__pe__lane19_strm0_data_valid ),      
               .std__pe__lane19_strm0_data_mask     ( std__pe__lane19_strm0_data_mask  ),      
               .pe__std__lane19_strm1_ready         ( pe__std__lane19_strm1_ready      ),      
               .std__pe__lane19_strm1_cntl          ( std__pe__lane19_strm1_cntl       ),      
               .std__pe__lane19_strm1_data          ( std__pe__lane19_strm1_data       ),      
               .std__pe__lane19_strm1_data_valid    ( std__pe__lane19_strm1_data_valid ),      
               .std__pe__lane19_strm1_data_mask     ( std__pe__lane19_strm1_data_mask  ),      
               // Lane 20                 
               .pe__std__lane20_strm0_ready         ( pe__std__lane20_strm0_ready      ),      
               .std__pe__lane20_strm0_cntl          ( std__pe__lane20_strm0_cntl       ),      
               .std__pe__lane20_strm0_data          ( std__pe__lane20_strm0_data       ),      
               .std__pe__lane20_strm0_data_valid    ( std__pe__lane20_strm0_data_valid ),      
               .std__pe__lane20_strm0_data_mask     ( std__pe__lane20_strm0_data_mask  ),      
               .pe__std__lane20_strm1_ready         ( pe__std__lane20_strm1_ready      ),      
               .std__pe__lane20_strm1_cntl          ( std__pe__lane20_strm1_cntl       ),      
               .std__pe__lane20_strm1_data          ( std__pe__lane20_strm1_data       ),      
               .std__pe__lane20_strm1_data_valid    ( std__pe__lane20_strm1_data_valid ),      
               .std__pe__lane20_strm1_data_mask     ( std__pe__lane20_strm1_data_mask  ),      
               // Lane 21                 
               .pe__std__lane21_strm0_ready         ( pe__std__lane21_strm0_ready      ),      
               .std__pe__lane21_strm0_cntl          ( std__pe__lane21_strm0_cntl       ),      
               .std__pe__lane21_strm0_data          ( std__pe__lane21_strm0_data       ),      
               .std__pe__lane21_strm0_data_valid    ( std__pe__lane21_strm0_data_valid ),      
               .std__pe__lane21_strm0_data_mask     ( std__pe__lane21_strm0_data_mask  ),      
               .pe__std__lane21_strm1_ready         ( pe__std__lane21_strm1_ready      ),      
               .std__pe__lane21_strm1_cntl          ( std__pe__lane21_strm1_cntl       ),      
               .std__pe__lane21_strm1_data          ( std__pe__lane21_strm1_data       ),      
               .std__pe__lane21_strm1_data_valid    ( std__pe__lane21_strm1_data_valid ),      
               .std__pe__lane21_strm1_data_mask     ( std__pe__lane21_strm1_data_mask  ),      
               // Lane 22                 
               .pe__std__lane22_strm0_ready         ( pe__std__lane22_strm0_ready      ),      
               .std__pe__lane22_strm0_cntl          ( std__pe__lane22_strm0_cntl       ),      
               .std__pe__lane22_strm0_data          ( std__pe__lane22_strm0_data       ),      
               .std__pe__lane22_strm0_data_valid    ( std__pe__lane22_strm0_data_valid ),      
               .std__pe__lane22_strm0_data_mask     ( std__pe__lane22_strm0_data_mask  ),      
               .pe__std__lane22_strm1_ready         ( pe__std__lane22_strm1_ready      ),      
               .std__pe__lane22_strm1_cntl          ( std__pe__lane22_strm1_cntl       ),      
               .std__pe__lane22_strm1_data          ( std__pe__lane22_strm1_data       ),      
               .std__pe__lane22_strm1_data_valid    ( std__pe__lane22_strm1_data_valid ),      
               .std__pe__lane22_strm1_data_mask     ( std__pe__lane22_strm1_data_mask  ),      
               // Lane 23                 
               .pe__std__lane23_strm0_ready         ( pe__std__lane23_strm0_ready      ),      
               .std__pe__lane23_strm0_cntl          ( std__pe__lane23_strm0_cntl       ),      
               .std__pe__lane23_strm0_data          ( std__pe__lane23_strm0_data       ),      
               .std__pe__lane23_strm0_data_valid    ( std__pe__lane23_strm0_data_valid ),      
               .std__pe__lane23_strm0_data_mask     ( std__pe__lane23_strm0_data_mask  ),      
               .pe__std__lane23_strm1_ready         ( pe__std__lane23_strm1_ready      ),      
               .std__pe__lane23_strm1_cntl          ( std__pe__lane23_strm1_cntl       ),      
               .std__pe__lane23_strm1_data          ( std__pe__lane23_strm1_data       ),      
               .std__pe__lane23_strm1_data_valid    ( std__pe__lane23_strm1_data_valid ),      
               .std__pe__lane23_strm1_data_mask     ( std__pe__lane23_strm1_data_mask  ),      
               // Lane 24                 
               .pe__std__lane24_strm0_ready         ( pe__std__lane24_strm0_ready      ),      
               .std__pe__lane24_strm0_cntl          ( std__pe__lane24_strm0_cntl       ),      
               .std__pe__lane24_strm0_data          ( std__pe__lane24_strm0_data       ),      
               .std__pe__lane24_strm0_data_valid    ( std__pe__lane24_strm0_data_valid ),      
               .std__pe__lane24_strm0_data_mask     ( std__pe__lane24_strm0_data_mask  ),      
               .pe__std__lane24_strm1_ready         ( pe__std__lane24_strm1_ready      ),      
               .std__pe__lane24_strm1_cntl          ( std__pe__lane24_strm1_cntl       ),      
               .std__pe__lane24_strm1_data          ( std__pe__lane24_strm1_data       ),      
               .std__pe__lane24_strm1_data_valid    ( std__pe__lane24_strm1_data_valid ),      
               .std__pe__lane24_strm1_data_mask     ( std__pe__lane24_strm1_data_mask  ),      
               // Lane 25                 
               .pe__std__lane25_strm0_ready         ( pe__std__lane25_strm0_ready      ),      
               .std__pe__lane25_strm0_cntl          ( std__pe__lane25_strm0_cntl       ),      
               .std__pe__lane25_strm0_data          ( std__pe__lane25_strm0_data       ),      
               .std__pe__lane25_strm0_data_valid    ( std__pe__lane25_strm0_data_valid ),      
               .std__pe__lane25_strm0_data_mask     ( std__pe__lane25_strm0_data_mask  ),      
               .pe__std__lane25_strm1_ready         ( pe__std__lane25_strm1_ready      ),      
               .std__pe__lane25_strm1_cntl          ( std__pe__lane25_strm1_cntl       ),      
               .std__pe__lane25_strm1_data          ( std__pe__lane25_strm1_data       ),      
               .std__pe__lane25_strm1_data_valid    ( std__pe__lane25_strm1_data_valid ),      
               .std__pe__lane25_strm1_data_mask     ( std__pe__lane25_strm1_data_mask  ),      
               // Lane 26                 
               .pe__std__lane26_strm0_ready         ( pe__std__lane26_strm0_ready      ),      
               .std__pe__lane26_strm0_cntl          ( std__pe__lane26_strm0_cntl       ),      
               .std__pe__lane26_strm0_data          ( std__pe__lane26_strm0_data       ),      
               .std__pe__lane26_strm0_data_valid    ( std__pe__lane26_strm0_data_valid ),      
               .std__pe__lane26_strm0_data_mask     ( std__pe__lane26_strm0_data_mask  ),      
               .pe__std__lane26_strm1_ready         ( pe__std__lane26_strm1_ready      ),      
               .std__pe__lane26_strm1_cntl          ( std__pe__lane26_strm1_cntl       ),      
               .std__pe__lane26_strm1_data          ( std__pe__lane26_strm1_data       ),      
               .std__pe__lane26_strm1_data_valid    ( std__pe__lane26_strm1_data_valid ),      
               .std__pe__lane26_strm1_data_mask     ( std__pe__lane26_strm1_data_mask  ),      
               // Lane 27                 
               .pe__std__lane27_strm0_ready         ( pe__std__lane27_strm0_ready      ),      
               .std__pe__lane27_strm0_cntl          ( std__pe__lane27_strm0_cntl       ),      
               .std__pe__lane27_strm0_data          ( std__pe__lane27_strm0_data       ),      
               .std__pe__lane27_strm0_data_valid    ( std__pe__lane27_strm0_data_valid ),      
               .std__pe__lane27_strm0_data_mask     ( std__pe__lane27_strm0_data_mask  ),      
               .pe__std__lane27_strm1_ready         ( pe__std__lane27_strm1_ready      ),      
               .std__pe__lane27_strm1_cntl          ( std__pe__lane27_strm1_cntl       ),      
               .std__pe__lane27_strm1_data          ( std__pe__lane27_strm1_data       ),      
               .std__pe__lane27_strm1_data_valid    ( std__pe__lane27_strm1_data_valid ),      
               .std__pe__lane27_strm1_data_mask     ( std__pe__lane27_strm1_data_mask  ),      
               // Lane 28                 
               .pe__std__lane28_strm0_ready         ( pe__std__lane28_strm0_ready      ),      
               .std__pe__lane28_strm0_cntl          ( std__pe__lane28_strm0_cntl       ),      
               .std__pe__lane28_strm0_data          ( std__pe__lane28_strm0_data       ),      
               .std__pe__lane28_strm0_data_valid    ( std__pe__lane28_strm0_data_valid ),      
               .std__pe__lane28_strm0_data_mask     ( std__pe__lane28_strm0_data_mask  ),      
               .pe__std__lane28_strm1_ready         ( pe__std__lane28_strm1_ready      ),      
               .std__pe__lane28_strm1_cntl          ( std__pe__lane28_strm1_cntl       ),      
               .std__pe__lane28_strm1_data          ( std__pe__lane28_strm1_data       ),      
               .std__pe__lane28_strm1_data_valid    ( std__pe__lane28_strm1_data_valid ),      
               .std__pe__lane28_strm1_data_mask     ( std__pe__lane28_strm1_data_mask  ),      
               // Lane 29                 
               .pe__std__lane29_strm0_ready         ( pe__std__lane29_strm0_ready      ),      
               .std__pe__lane29_strm0_cntl          ( std__pe__lane29_strm0_cntl       ),      
               .std__pe__lane29_strm0_data          ( std__pe__lane29_strm0_data       ),      
               .std__pe__lane29_strm0_data_valid    ( std__pe__lane29_strm0_data_valid ),      
               .std__pe__lane29_strm0_data_mask     ( std__pe__lane29_strm0_data_mask  ),      
               .pe__std__lane29_strm1_ready         ( pe__std__lane29_strm1_ready      ),      
               .std__pe__lane29_strm1_cntl          ( std__pe__lane29_strm1_cntl       ),      
               .std__pe__lane29_strm1_data          ( std__pe__lane29_strm1_data       ),      
               .std__pe__lane29_strm1_data_valid    ( std__pe__lane29_strm1_data_valid ),      
               .std__pe__lane29_strm1_data_mask     ( std__pe__lane29_strm1_data_mask  ),      
               // Lane 30                 
               .pe__std__lane30_strm0_ready         ( pe__std__lane30_strm0_ready      ),      
               .std__pe__lane30_strm0_cntl          ( std__pe__lane30_strm0_cntl       ),      
               .std__pe__lane30_strm0_data          ( std__pe__lane30_strm0_data       ),      
               .std__pe__lane30_strm0_data_valid    ( std__pe__lane30_strm0_data_valid ),      
               .std__pe__lane30_strm0_data_mask     ( std__pe__lane30_strm0_data_mask  ),      
               .pe__std__lane30_strm1_ready         ( pe__std__lane30_strm1_ready      ),      
               .std__pe__lane30_strm1_cntl          ( std__pe__lane30_strm1_cntl       ),      
               .std__pe__lane30_strm1_data          ( std__pe__lane30_strm1_data       ),      
               .std__pe__lane30_strm1_data_valid    ( std__pe__lane30_strm1_data_valid ),      
               .std__pe__lane30_strm1_data_mask     ( std__pe__lane30_strm1_data_mask  ),      
               // Lane 31                 
               .pe__std__lane31_strm0_ready         ( pe__std__lane31_strm0_ready      ),      
               .std__pe__lane31_strm0_cntl          ( std__pe__lane31_strm0_cntl       ),      
               .std__pe__lane31_strm0_data          ( std__pe__lane31_strm0_data       ),      
               .std__pe__lane31_strm0_data_valid    ( std__pe__lane31_strm0_data_valid ),      
               .std__pe__lane31_strm0_data_mask     ( std__pe__lane31_strm0_data_mask  ),      
               .pe__std__lane31_strm1_ready         ( pe__std__lane31_strm1_ready      ),      
               .std__pe__lane31_strm1_cntl          ( std__pe__lane31_strm1_cntl       ),      
               .std__pe__lane31_strm1_data          ( std__pe__lane31_strm1_data       ),      
               .std__pe__lane31_strm1_data_valid    ( std__pe__lane31_strm1_data_valid ),      
               .std__pe__lane31_strm1_data_mask     ( std__pe__lane31_strm1_data_mask  ),      