
        begin
          forever
            begin
              // Observe NoC packets received by manager 0
              @(vLocalFromNoC[0].cb_p);
              if ((vLocalFromNoC[0].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[0].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [0] = new();
                  local_noc_pkt_rcvd [0].header_destination_address  = vLocalFromNoC[0].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [0].header_source               = vLocalFromNoC[0].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [0].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 0, vLocalFromNoC[0].noc__locl__dp_mgrId);
                  noc2mgr_p [0].put(local_noc_pkt_rcvd [0]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 1
              @(vLocalFromNoC[1].cb_p);
              if ((vLocalFromNoC[1].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[1].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [1] = new();
                  local_noc_pkt_rcvd [1].header_destination_address  = vLocalFromNoC[1].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [1].header_source               = vLocalFromNoC[1].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [1].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 1, vLocalFromNoC[1].noc__locl__dp_mgrId);
                  noc2mgr_p [1].put(local_noc_pkt_rcvd [1]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 2
              @(vLocalFromNoC[2].cb_p);
              if ((vLocalFromNoC[2].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[2].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [2] = new();
                  local_noc_pkt_rcvd [2].header_destination_address  = vLocalFromNoC[2].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [2].header_source               = vLocalFromNoC[2].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [2].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 2, vLocalFromNoC[2].noc__locl__dp_mgrId);
                  noc2mgr_p [2].put(local_noc_pkt_rcvd [2]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 3
              @(vLocalFromNoC[3].cb_p);
              if ((vLocalFromNoC[3].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[3].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [3] = new();
                  local_noc_pkt_rcvd [3].header_destination_address  = vLocalFromNoC[3].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [3].header_source               = vLocalFromNoC[3].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [3].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 3, vLocalFromNoC[3].noc__locl__dp_mgrId);
                  noc2mgr_p [3].put(local_noc_pkt_rcvd [3]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 4
              @(vLocalFromNoC[4].cb_p);
              if ((vLocalFromNoC[4].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[4].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [4] = new();
                  local_noc_pkt_rcvd [4].header_destination_address  = vLocalFromNoC[4].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [4].header_source               = vLocalFromNoC[4].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [4].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 4, vLocalFromNoC[4].noc__locl__dp_mgrId);
                  noc2mgr_p [4].put(local_noc_pkt_rcvd [4]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 5
              @(vLocalFromNoC[5].cb_p);
              if ((vLocalFromNoC[5].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[5].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [5] = new();
                  local_noc_pkt_rcvd [5].header_destination_address  = vLocalFromNoC[5].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [5].header_source               = vLocalFromNoC[5].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [5].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 5, vLocalFromNoC[5].noc__locl__dp_mgrId);
                  noc2mgr_p [5].put(local_noc_pkt_rcvd [5]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 6
              @(vLocalFromNoC[6].cb_p);
              if ((vLocalFromNoC[6].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[6].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [6] = new();
                  local_noc_pkt_rcvd [6].header_destination_address  = vLocalFromNoC[6].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [6].header_source               = vLocalFromNoC[6].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [6].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 6, vLocalFromNoC[6].noc__locl__dp_mgrId);
                  noc2mgr_p [6].put(local_noc_pkt_rcvd [6]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 7
              @(vLocalFromNoC[7].cb_p);
              if ((vLocalFromNoC[7].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[7].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [7] = new();
                  local_noc_pkt_rcvd [7].header_destination_address  = vLocalFromNoC[7].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [7].header_source               = vLocalFromNoC[7].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [7].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 7, vLocalFromNoC[7].noc__locl__dp_mgrId);
                  noc2mgr_p [7].put(local_noc_pkt_rcvd [7]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 8
              @(vLocalFromNoC[8].cb_p);
              if ((vLocalFromNoC[8].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[8].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [8] = new();
                  local_noc_pkt_rcvd [8].header_destination_address  = vLocalFromNoC[8].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [8].header_source               = vLocalFromNoC[8].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [8].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 8, vLocalFromNoC[8].noc__locl__dp_mgrId);
                  noc2mgr_p [8].put(local_noc_pkt_rcvd [8]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 9
              @(vLocalFromNoC[9].cb_p);
              if ((vLocalFromNoC[9].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[9].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [9] = new();
                  local_noc_pkt_rcvd [9].header_destination_address  = vLocalFromNoC[9].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [9].header_source               = vLocalFromNoC[9].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [9].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 9, vLocalFromNoC[9].noc__locl__dp_mgrId);
                  noc2mgr_p [9].put(local_noc_pkt_rcvd [9]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 10
              @(vLocalFromNoC[10].cb_p);
              if ((vLocalFromNoC[10].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[10].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [10] = new();
                  local_noc_pkt_rcvd [10].header_destination_address  = vLocalFromNoC[10].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [10].header_source               = vLocalFromNoC[10].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [10].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 10, vLocalFromNoC[10].noc__locl__dp_mgrId);
                  noc2mgr_p [10].put(local_noc_pkt_rcvd [10]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 11
              @(vLocalFromNoC[11].cb_p);
              if ((vLocalFromNoC[11].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[11].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [11] = new();
                  local_noc_pkt_rcvd [11].header_destination_address  = vLocalFromNoC[11].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [11].header_source               = vLocalFromNoC[11].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [11].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 11, vLocalFromNoC[11].noc__locl__dp_mgrId);
                  noc2mgr_p [11].put(local_noc_pkt_rcvd [11]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 12
              @(vLocalFromNoC[12].cb_p);
              if ((vLocalFromNoC[12].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[12].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [12] = new();
                  local_noc_pkt_rcvd [12].header_destination_address  = vLocalFromNoC[12].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [12].header_source               = vLocalFromNoC[12].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [12].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 12, vLocalFromNoC[12].noc__locl__dp_mgrId);
                  noc2mgr_p [12].put(local_noc_pkt_rcvd [12]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 13
              @(vLocalFromNoC[13].cb_p);
              if ((vLocalFromNoC[13].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[13].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [13] = new();
                  local_noc_pkt_rcvd [13].header_destination_address  = vLocalFromNoC[13].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [13].header_source               = vLocalFromNoC[13].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [13].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 13, vLocalFromNoC[13].noc__locl__dp_mgrId);
                  noc2mgr_p [13].put(local_noc_pkt_rcvd [13]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 14
              @(vLocalFromNoC[14].cb_p);
              if ((vLocalFromNoC[14].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[14].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [14] = new();
                  local_noc_pkt_rcvd [14].header_destination_address  = vLocalFromNoC[14].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [14].header_source               = vLocalFromNoC[14].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [14].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 14, vLocalFromNoC[14].noc__locl__dp_mgrId);
                  noc2mgr_p [14].put(local_noc_pkt_rcvd [14]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 15
              @(vLocalFromNoC[15].cb_p);
              if ((vLocalFromNoC[15].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[15].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [15] = new();
                  local_noc_pkt_rcvd [15].header_destination_address  = vLocalFromNoC[15].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [15].header_source               = vLocalFromNoC[15].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [15].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 15, vLocalFromNoC[15].noc__locl__dp_mgrId);
                  noc2mgr_p [15].put(local_noc_pkt_rcvd [15]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 16
              @(vLocalFromNoC[16].cb_p);
              if ((vLocalFromNoC[16].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[16].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [16] = new();
                  local_noc_pkt_rcvd [16].header_destination_address  = vLocalFromNoC[16].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [16].header_source               = vLocalFromNoC[16].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [16].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 16, vLocalFromNoC[16].noc__locl__dp_mgrId);
                  noc2mgr_p [16].put(local_noc_pkt_rcvd [16]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 17
              @(vLocalFromNoC[17].cb_p);
              if ((vLocalFromNoC[17].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[17].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [17] = new();
                  local_noc_pkt_rcvd [17].header_destination_address  = vLocalFromNoC[17].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [17].header_source               = vLocalFromNoC[17].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [17].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 17, vLocalFromNoC[17].noc__locl__dp_mgrId);
                  noc2mgr_p [17].put(local_noc_pkt_rcvd [17]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 18
              @(vLocalFromNoC[18].cb_p);
              if ((vLocalFromNoC[18].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[18].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [18] = new();
                  local_noc_pkt_rcvd [18].header_destination_address  = vLocalFromNoC[18].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [18].header_source               = vLocalFromNoC[18].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [18].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 18, vLocalFromNoC[18].noc__locl__dp_mgrId);
                  noc2mgr_p [18].put(local_noc_pkt_rcvd [18]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 19
              @(vLocalFromNoC[19].cb_p);
              if ((vLocalFromNoC[19].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[19].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [19] = new();
                  local_noc_pkt_rcvd [19].header_destination_address  = vLocalFromNoC[19].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [19].header_source               = vLocalFromNoC[19].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [19].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 19, vLocalFromNoC[19].noc__locl__dp_mgrId);
                  noc2mgr_p [19].put(local_noc_pkt_rcvd [19]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 20
              @(vLocalFromNoC[20].cb_p);
              if ((vLocalFromNoC[20].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[20].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [20] = new();
                  local_noc_pkt_rcvd [20].header_destination_address  = vLocalFromNoC[20].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [20].header_source               = vLocalFromNoC[20].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [20].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 20, vLocalFromNoC[20].noc__locl__dp_mgrId);
                  noc2mgr_p [20].put(local_noc_pkt_rcvd [20]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 21
              @(vLocalFromNoC[21].cb_p);
              if ((vLocalFromNoC[21].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[21].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [21] = new();
                  local_noc_pkt_rcvd [21].header_destination_address  = vLocalFromNoC[21].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [21].header_source               = vLocalFromNoC[21].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [21].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 21, vLocalFromNoC[21].noc__locl__dp_mgrId);
                  noc2mgr_p [21].put(local_noc_pkt_rcvd [21]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 22
              @(vLocalFromNoC[22].cb_p);
              if ((vLocalFromNoC[22].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[22].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [22] = new();
                  local_noc_pkt_rcvd [22].header_destination_address  = vLocalFromNoC[22].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [22].header_source               = vLocalFromNoC[22].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [22].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 22, vLocalFromNoC[22].noc__locl__dp_mgrId);
                  noc2mgr_p [22].put(local_noc_pkt_rcvd [22]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 23
              @(vLocalFromNoC[23].cb_p);
              if ((vLocalFromNoC[23].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[23].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [23] = new();
                  local_noc_pkt_rcvd [23].header_destination_address  = vLocalFromNoC[23].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [23].header_source               = vLocalFromNoC[23].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [23].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 23, vLocalFromNoC[23].noc__locl__dp_mgrId);
                  noc2mgr_p [23].put(local_noc_pkt_rcvd [23]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 24
              @(vLocalFromNoC[24].cb_p);
              if ((vLocalFromNoC[24].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[24].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [24] = new();
                  local_noc_pkt_rcvd [24].header_destination_address  = vLocalFromNoC[24].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [24].header_source               = vLocalFromNoC[24].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [24].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 24, vLocalFromNoC[24].noc__locl__dp_mgrId);
                  noc2mgr_p [24].put(local_noc_pkt_rcvd [24]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 25
              @(vLocalFromNoC[25].cb_p);
              if ((vLocalFromNoC[25].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[25].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [25] = new();
                  local_noc_pkt_rcvd [25].header_destination_address  = vLocalFromNoC[25].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [25].header_source               = vLocalFromNoC[25].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [25].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 25, vLocalFromNoC[25].noc__locl__dp_mgrId);
                  noc2mgr_p [25].put(local_noc_pkt_rcvd [25]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 26
              @(vLocalFromNoC[26].cb_p);
              if ((vLocalFromNoC[26].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[26].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [26] = new();
                  local_noc_pkt_rcvd [26].header_destination_address  = vLocalFromNoC[26].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [26].header_source               = vLocalFromNoC[26].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [26].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 26, vLocalFromNoC[26].noc__locl__dp_mgrId);
                  noc2mgr_p [26].put(local_noc_pkt_rcvd [26]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 27
              @(vLocalFromNoC[27].cb_p);
              if ((vLocalFromNoC[27].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[27].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [27] = new();
                  local_noc_pkt_rcvd [27].header_destination_address  = vLocalFromNoC[27].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [27].header_source               = vLocalFromNoC[27].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [27].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 27, vLocalFromNoC[27].noc__locl__dp_mgrId);
                  noc2mgr_p [27].put(local_noc_pkt_rcvd [27]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 28
              @(vLocalFromNoC[28].cb_p);
              if ((vLocalFromNoC[28].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[28].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [28] = new();
                  local_noc_pkt_rcvd [28].header_destination_address  = vLocalFromNoC[28].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [28].header_source               = vLocalFromNoC[28].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [28].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 28, vLocalFromNoC[28].noc__locl__dp_mgrId);
                  noc2mgr_p [28].put(local_noc_pkt_rcvd [28]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 29
              @(vLocalFromNoC[29].cb_p);
              if ((vLocalFromNoC[29].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[29].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [29] = new();
                  local_noc_pkt_rcvd [29].header_destination_address  = vLocalFromNoC[29].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [29].header_source               = vLocalFromNoC[29].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [29].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 29, vLocalFromNoC[29].noc__locl__dp_mgrId);
                  noc2mgr_p [29].put(local_noc_pkt_rcvd [29]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 30
              @(vLocalFromNoC[30].cb_p);
              if ((vLocalFromNoC[30].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[30].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [30] = new();
                  local_noc_pkt_rcvd [30].header_destination_address  = vLocalFromNoC[30].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [30].header_source               = vLocalFromNoC[30].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [30].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 30, vLocalFromNoC[30].noc__locl__dp_mgrId);
                  noc2mgr_p [30].put(local_noc_pkt_rcvd [30]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 31
              @(vLocalFromNoC[31].cb_p);
              if ((vLocalFromNoC[31].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[31].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [31] = new();
                  local_noc_pkt_rcvd [31].header_destination_address  = vLocalFromNoC[31].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [31].header_source               = vLocalFromNoC[31].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [31].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 31, vLocalFromNoC[31].noc__locl__dp_mgrId);
                  noc2mgr_p [31].put(local_noc_pkt_rcvd [31]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 32
              @(vLocalFromNoC[32].cb_p);
              if ((vLocalFromNoC[32].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[32].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [32] = new();
                  local_noc_pkt_rcvd [32].header_destination_address  = vLocalFromNoC[32].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [32].header_source               = vLocalFromNoC[32].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [32].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 32, vLocalFromNoC[32].noc__locl__dp_mgrId);
                  noc2mgr_p [32].put(local_noc_pkt_rcvd [32]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 33
              @(vLocalFromNoC[33].cb_p);
              if ((vLocalFromNoC[33].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[33].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [33] = new();
                  local_noc_pkt_rcvd [33].header_destination_address  = vLocalFromNoC[33].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [33].header_source               = vLocalFromNoC[33].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [33].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 33, vLocalFromNoC[33].noc__locl__dp_mgrId);
                  noc2mgr_p [33].put(local_noc_pkt_rcvd [33]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 34
              @(vLocalFromNoC[34].cb_p);
              if ((vLocalFromNoC[34].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[34].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [34] = new();
                  local_noc_pkt_rcvd [34].header_destination_address  = vLocalFromNoC[34].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [34].header_source               = vLocalFromNoC[34].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [34].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 34, vLocalFromNoC[34].noc__locl__dp_mgrId);
                  noc2mgr_p [34].put(local_noc_pkt_rcvd [34]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 35
              @(vLocalFromNoC[35].cb_p);
              if ((vLocalFromNoC[35].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[35].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [35] = new();
                  local_noc_pkt_rcvd [35].header_destination_address  = vLocalFromNoC[35].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [35].header_source               = vLocalFromNoC[35].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [35].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 35, vLocalFromNoC[35].noc__locl__dp_mgrId);
                  noc2mgr_p [35].put(local_noc_pkt_rcvd [35]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 36
              @(vLocalFromNoC[36].cb_p);
              if ((vLocalFromNoC[36].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[36].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [36] = new();
                  local_noc_pkt_rcvd [36].header_destination_address  = vLocalFromNoC[36].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [36].header_source               = vLocalFromNoC[36].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [36].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 36, vLocalFromNoC[36].noc__locl__dp_mgrId);
                  noc2mgr_p [36].put(local_noc_pkt_rcvd [36]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 37
              @(vLocalFromNoC[37].cb_p);
              if ((vLocalFromNoC[37].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[37].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [37] = new();
                  local_noc_pkt_rcvd [37].header_destination_address  = vLocalFromNoC[37].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [37].header_source               = vLocalFromNoC[37].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [37].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 37, vLocalFromNoC[37].noc__locl__dp_mgrId);
                  noc2mgr_p [37].put(local_noc_pkt_rcvd [37]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 38
              @(vLocalFromNoC[38].cb_p);
              if ((vLocalFromNoC[38].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[38].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [38] = new();
                  local_noc_pkt_rcvd [38].header_destination_address  = vLocalFromNoC[38].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [38].header_source               = vLocalFromNoC[38].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [38].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 38, vLocalFromNoC[38].noc__locl__dp_mgrId);
                  noc2mgr_p [38].put(local_noc_pkt_rcvd [38]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 39
              @(vLocalFromNoC[39].cb_p);
              if ((vLocalFromNoC[39].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[39].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [39] = new();
                  local_noc_pkt_rcvd [39].header_destination_address  = vLocalFromNoC[39].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [39].header_source               = vLocalFromNoC[39].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [39].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 39, vLocalFromNoC[39].noc__locl__dp_mgrId);
                  noc2mgr_p [39].put(local_noc_pkt_rcvd [39]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 40
              @(vLocalFromNoC[40].cb_p);
              if ((vLocalFromNoC[40].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[40].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [40] = new();
                  local_noc_pkt_rcvd [40].header_destination_address  = vLocalFromNoC[40].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [40].header_source               = vLocalFromNoC[40].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [40].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 40, vLocalFromNoC[40].noc__locl__dp_mgrId);
                  noc2mgr_p [40].put(local_noc_pkt_rcvd [40]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 41
              @(vLocalFromNoC[41].cb_p);
              if ((vLocalFromNoC[41].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[41].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [41] = new();
                  local_noc_pkt_rcvd [41].header_destination_address  = vLocalFromNoC[41].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [41].header_source               = vLocalFromNoC[41].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [41].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 41, vLocalFromNoC[41].noc__locl__dp_mgrId);
                  noc2mgr_p [41].put(local_noc_pkt_rcvd [41]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 42
              @(vLocalFromNoC[42].cb_p);
              if ((vLocalFromNoC[42].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[42].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [42] = new();
                  local_noc_pkt_rcvd [42].header_destination_address  = vLocalFromNoC[42].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [42].header_source               = vLocalFromNoC[42].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [42].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 42, vLocalFromNoC[42].noc__locl__dp_mgrId);
                  noc2mgr_p [42].put(local_noc_pkt_rcvd [42]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 43
              @(vLocalFromNoC[43].cb_p);
              if ((vLocalFromNoC[43].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[43].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [43] = new();
                  local_noc_pkt_rcvd [43].header_destination_address  = vLocalFromNoC[43].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [43].header_source               = vLocalFromNoC[43].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [43].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 43, vLocalFromNoC[43].noc__locl__dp_mgrId);
                  noc2mgr_p [43].put(local_noc_pkt_rcvd [43]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 44
              @(vLocalFromNoC[44].cb_p);
              if ((vLocalFromNoC[44].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[44].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [44] = new();
                  local_noc_pkt_rcvd [44].header_destination_address  = vLocalFromNoC[44].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [44].header_source               = vLocalFromNoC[44].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [44].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 44, vLocalFromNoC[44].noc__locl__dp_mgrId);
                  noc2mgr_p [44].put(local_noc_pkt_rcvd [44]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 45
              @(vLocalFromNoC[45].cb_p);
              if ((vLocalFromNoC[45].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[45].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [45] = new();
                  local_noc_pkt_rcvd [45].header_destination_address  = vLocalFromNoC[45].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [45].header_source               = vLocalFromNoC[45].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [45].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 45, vLocalFromNoC[45].noc__locl__dp_mgrId);
                  noc2mgr_p [45].put(local_noc_pkt_rcvd [45]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 46
              @(vLocalFromNoC[46].cb_p);
              if ((vLocalFromNoC[46].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[46].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [46] = new();
                  local_noc_pkt_rcvd [46].header_destination_address  = vLocalFromNoC[46].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [46].header_source               = vLocalFromNoC[46].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [46].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 46, vLocalFromNoC[46].noc__locl__dp_mgrId);
                  noc2mgr_p [46].put(local_noc_pkt_rcvd [46]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 47
              @(vLocalFromNoC[47].cb_p);
              if ((vLocalFromNoC[47].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[47].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [47] = new();
                  local_noc_pkt_rcvd [47].header_destination_address  = vLocalFromNoC[47].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [47].header_source               = vLocalFromNoC[47].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [47].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 47, vLocalFromNoC[47].noc__locl__dp_mgrId);
                  noc2mgr_p [47].put(local_noc_pkt_rcvd [47]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 48
              @(vLocalFromNoC[48].cb_p);
              if ((vLocalFromNoC[48].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[48].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [48] = new();
                  local_noc_pkt_rcvd [48].header_destination_address  = vLocalFromNoC[48].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [48].header_source               = vLocalFromNoC[48].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [48].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 48, vLocalFromNoC[48].noc__locl__dp_mgrId);
                  noc2mgr_p [48].put(local_noc_pkt_rcvd [48]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 49
              @(vLocalFromNoC[49].cb_p);
              if ((vLocalFromNoC[49].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[49].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [49] = new();
                  local_noc_pkt_rcvd [49].header_destination_address  = vLocalFromNoC[49].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [49].header_source               = vLocalFromNoC[49].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [49].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 49, vLocalFromNoC[49].noc__locl__dp_mgrId);
                  noc2mgr_p [49].put(local_noc_pkt_rcvd [49]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 50
              @(vLocalFromNoC[50].cb_p);
              if ((vLocalFromNoC[50].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[50].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [50] = new();
                  local_noc_pkt_rcvd [50].header_destination_address  = vLocalFromNoC[50].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [50].header_source               = vLocalFromNoC[50].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [50].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 50, vLocalFromNoC[50].noc__locl__dp_mgrId);
                  noc2mgr_p [50].put(local_noc_pkt_rcvd [50]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 51
              @(vLocalFromNoC[51].cb_p);
              if ((vLocalFromNoC[51].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[51].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [51] = new();
                  local_noc_pkt_rcvd [51].header_destination_address  = vLocalFromNoC[51].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [51].header_source               = vLocalFromNoC[51].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [51].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 51, vLocalFromNoC[51].noc__locl__dp_mgrId);
                  noc2mgr_p [51].put(local_noc_pkt_rcvd [51]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 52
              @(vLocalFromNoC[52].cb_p);
              if ((vLocalFromNoC[52].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[52].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [52] = new();
                  local_noc_pkt_rcvd [52].header_destination_address  = vLocalFromNoC[52].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [52].header_source               = vLocalFromNoC[52].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [52].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 52, vLocalFromNoC[52].noc__locl__dp_mgrId);
                  noc2mgr_p [52].put(local_noc_pkt_rcvd [52]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 53
              @(vLocalFromNoC[53].cb_p);
              if ((vLocalFromNoC[53].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[53].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [53] = new();
                  local_noc_pkt_rcvd [53].header_destination_address  = vLocalFromNoC[53].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [53].header_source               = vLocalFromNoC[53].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [53].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 53, vLocalFromNoC[53].noc__locl__dp_mgrId);
                  noc2mgr_p [53].put(local_noc_pkt_rcvd [53]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 54
              @(vLocalFromNoC[54].cb_p);
              if ((vLocalFromNoC[54].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[54].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [54] = new();
                  local_noc_pkt_rcvd [54].header_destination_address  = vLocalFromNoC[54].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [54].header_source               = vLocalFromNoC[54].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [54].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 54, vLocalFromNoC[54].noc__locl__dp_mgrId);
                  noc2mgr_p [54].put(local_noc_pkt_rcvd [54]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 55
              @(vLocalFromNoC[55].cb_p);
              if ((vLocalFromNoC[55].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[55].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [55] = new();
                  local_noc_pkt_rcvd [55].header_destination_address  = vLocalFromNoC[55].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [55].header_source               = vLocalFromNoC[55].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [55].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 55, vLocalFromNoC[55].noc__locl__dp_mgrId);
                  noc2mgr_p [55].put(local_noc_pkt_rcvd [55]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 56
              @(vLocalFromNoC[56].cb_p);
              if ((vLocalFromNoC[56].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[56].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [56] = new();
                  local_noc_pkt_rcvd [56].header_destination_address  = vLocalFromNoC[56].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [56].header_source               = vLocalFromNoC[56].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [56].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 56, vLocalFromNoC[56].noc__locl__dp_mgrId);
                  noc2mgr_p [56].put(local_noc_pkt_rcvd [56]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 57
              @(vLocalFromNoC[57].cb_p);
              if ((vLocalFromNoC[57].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[57].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [57] = new();
                  local_noc_pkt_rcvd [57].header_destination_address  = vLocalFromNoC[57].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [57].header_source               = vLocalFromNoC[57].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [57].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 57, vLocalFromNoC[57].noc__locl__dp_mgrId);
                  noc2mgr_p [57].put(local_noc_pkt_rcvd [57]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 58
              @(vLocalFromNoC[58].cb_p);
              if ((vLocalFromNoC[58].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[58].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [58] = new();
                  local_noc_pkt_rcvd [58].header_destination_address  = vLocalFromNoC[58].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [58].header_source               = vLocalFromNoC[58].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [58].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 58, vLocalFromNoC[58].noc__locl__dp_mgrId);
                  noc2mgr_p [58].put(local_noc_pkt_rcvd [58]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 59
              @(vLocalFromNoC[59].cb_p);
              if ((vLocalFromNoC[59].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[59].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [59] = new();
                  local_noc_pkt_rcvd [59].header_destination_address  = vLocalFromNoC[59].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [59].header_source               = vLocalFromNoC[59].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [59].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 59, vLocalFromNoC[59].noc__locl__dp_mgrId);
                  noc2mgr_p [59].put(local_noc_pkt_rcvd [59]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 60
              @(vLocalFromNoC[60].cb_p);
              if ((vLocalFromNoC[60].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[60].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [60] = new();
                  local_noc_pkt_rcvd [60].header_destination_address  = vLocalFromNoC[60].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [60].header_source               = vLocalFromNoC[60].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [60].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 60, vLocalFromNoC[60].noc__locl__dp_mgrId);
                  noc2mgr_p [60].put(local_noc_pkt_rcvd [60]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 61
              @(vLocalFromNoC[61].cb_p);
              if ((vLocalFromNoC[61].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[61].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [61] = new();
                  local_noc_pkt_rcvd [61].header_destination_address  = vLocalFromNoC[61].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [61].header_source               = vLocalFromNoC[61].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [61].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 61, vLocalFromNoC[61].noc__locl__dp_mgrId);
                  noc2mgr_p [61].put(local_noc_pkt_rcvd [61]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 62
              @(vLocalFromNoC[62].cb_p);
              if ((vLocalFromNoC[62].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[62].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [62] = new();
                  local_noc_pkt_rcvd [62].header_destination_address  = vLocalFromNoC[62].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [62].header_source               = vLocalFromNoC[62].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [62].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 62, vLocalFromNoC[62].noc__locl__dp_mgrId);
                  noc2mgr_p [62].put(local_noc_pkt_rcvd [62]);
                end
            end
        end
    
        begin
          forever
            begin
              // Observe NoC packets received by manager 63
              @(vLocalFromNoC[63].cb_p);
              if ((vLocalFromNoC[63].noc__locl__dp_valid == 1'b1) && (vLocalFromNoC[63].noc__locl__dp_cntl == 2'b01))
                begin
                  local_noc_pkt_rcvd [63] = new();
                  local_noc_pkt_rcvd [63].header_destination_address  = vLocalFromNoC[63].noc__locl__dp_data     ;
                  local_noc_pkt_rcvd [63].header_source               = vLocalFromNoC[63].noc__locl__dp_mgrId    ;
                  local_noc_pkt_rcvd [63].header_priority             = 1'b1                                   ;  // _dp is hi-priority
                  $display ("@%0t::%s:%0d:: INFO: Packet being received by {%0d} from {%0d}", $time, `__FILE__, `__LINE__, 63, vLocalFromNoC[63].noc__locl__dp_mgrId);
                  noc2mgr_p [63].put(local_noc_pkt_rcvd [63]);
                end
            end
        end
    