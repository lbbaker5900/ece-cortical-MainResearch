
  // General control and status                                                   
  input                                         mgr0__sys__allSynchronized     ;
  output                                        sys__mgr0__thisSynchronized    ;
  output                                        sys__mgr0__ready               ;
  output                                        sys__mgr0__complete            ;

  output                                        sys__pe0__allSynchronized     ;
  input                                         pe0__sys__thisSynchronized    ;
  input                                         pe0__sys__ready               ;
  input                                         pe0__sys__complete            ;

  // General control and status                                                   
  input                                         mgr1__sys__allSynchronized     ;
  output                                        sys__mgr1__thisSynchronized    ;
  output                                        sys__mgr1__ready               ;
  output                                        sys__mgr1__complete            ;

  output                                        sys__pe1__allSynchronized     ;
  input                                         pe1__sys__thisSynchronized    ;
  input                                         pe1__sys__ready               ;
  input                                         pe1__sys__complete            ;

  // General control and status                                                   
  input                                         mgr2__sys__allSynchronized     ;
  output                                        sys__mgr2__thisSynchronized    ;
  output                                        sys__mgr2__ready               ;
  output                                        sys__mgr2__complete            ;

  output                                        sys__pe2__allSynchronized     ;
  input                                         pe2__sys__thisSynchronized    ;
  input                                         pe2__sys__ready               ;
  input                                         pe2__sys__complete            ;

  // General control and status                                                   
  input                                         mgr3__sys__allSynchronized     ;
  output                                        sys__mgr3__thisSynchronized    ;
  output                                        sys__mgr3__ready               ;
  output                                        sys__mgr3__complete            ;

  output                                        sys__pe3__allSynchronized     ;
  input                                         pe3__sys__thisSynchronized    ;
  input                                         pe3__sys__ready               ;
  input                                         pe3__sys__complete            ;

  // General control and status                                                   
  input                                         mgr4__sys__allSynchronized     ;
  output                                        sys__mgr4__thisSynchronized    ;
  output                                        sys__mgr4__ready               ;
  output                                        sys__mgr4__complete            ;

  output                                        sys__pe4__allSynchronized     ;
  input                                         pe4__sys__thisSynchronized    ;
  input                                         pe4__sys__ready               ;
  input                                         pe4__sys__complete            ;

  // General control and status                                                   
  input                                         mgr5__sys__allSynchronized     ;
  output                                        sys__mgr5__thisSynchronized    ;
  output                                        sys__mgr5__ready               ;
  output                                        sys__mgr5__complete            ;

  output                                        sys__pe5__allSynchronized     ;
  input                                         pe5__sys__thisSynchronized    ;
  input                                         pe5__sys__ready               ;
  input                                         pe5__sys__complete            ;

  // General control and status                                                   
  input                                         mgr6__sys__allSynchronized     ;
  output                                        sys__mgr6__thisSynchronized    ;
  output                                        sys__mgr6__ready               ;
  output                                        sys__mgr6__complete            ;

  output                                        sys__pe6__allSynchronized     ;
  input                                         pe6__sys__thisSynchronized    ;
  input                                         pe6__sys__ready               ;
  input                                         pe6__sys__complete            ;

  // General control and status                                                   
  input                                         mgr7__sys__allSynchronized     ;
  output                                        sys__mgr7__thisSynchronized    ;
  output                                        sys__mgr7__ready               ;
  output                                        sys__mgr7__complete            ;

  output                                        sys__pe7__allSynchronized     ;
  input                                         pe7__sys__thisSynchronized    ;
  input                                         pe7__sys__ready               ;
  input                                         pe7__sys__complete            ;

  // General control and status                                                   
  input                                         mgr8__sys__allSynchronized     ;
  output                                        sys__mgr8__thisSynchronized    ;
  output                                        sys__mgr8__ready               ;
  output                                        sys__mgr8__complete            ;

  output                                        sys__pe8__allSynchronized     ;
  input                                         pe8__sys__thisSynchronized    ;
  input                                         pe8__sys__ready               ;
  input                                         pe8__sys__complete            ;

  // General control and status                                                   
  input                                         mgr9__sys__allSynchronized     ;
  output                                        sys__mgr9__thisSynchronized    ;
  output                                        sys__mgr9__ready               ;
  output                                        sys__mgr9__complete            ;

  output                                        sys__pe9__allSynchronized     ;
  input                                         pe9__sys__thisSynchronized    ;
  input                                         pe9__sys__ready               ;
  input                                         pe9__sys__complete            ;

  // General control and status                                                   
  input                                         mgr10__sys__allSynchronized     ;
  output                                        sys__mgr10__thisSynchronized    ;
  output                                        sys__mgr10__ready               ;
  output                                        sys__mgr10__complete            ;

  output                                        sys__pe10__allSynchronized     ;
  input                                         pe10__sys__thisSynchronized    ;
  input                                         pe10__sys__ready               ;
  input                                         pe10__sys__complete            ;

  // General control and status                                                   
  input                                         mgr11__sys__allSynchronized     ;
  output                                        sys__mgr11__thisSynchronized    ;
  output                                        sys__mgr11__ready               ;
  output                                        sys__mgr11__complete            ;

  output                                        sys__pe11__allSynchronized     ;
  input                                         pe11__sys__thisSynchronized    ;
  input                                         pe11__sys__ready               ;
  input                                         pe11__sys__complete            ;

  // General control and status                                                   
  input                                         mgr12__sys__allSynchronized     ;
  output                                        sys__mgr12__thisSynchronized    ;
  output                                        sys__mgr12__ready               ;
  output                                        sys__mgr12__complete            ;

  output                                        sys__pe12__allSynchronized     ;
  input                                         pe12__sys__thisSynchronized    ;
  input                                         pe12__sys__ready               ;
  input                                         pe12__sys__complete            ;

  // General control and status                                                   
  input                                         mgr13__sys__allSynchronized     ;
  output                                        sys__mgr13__thisSynchronized    ;
  output                                        sys__mgr13__ready               ;
  output                                        sys__mgr13__complete            ;

  output                                        sys__pe13__allSynchronized     ;
  input                                         pe13__sys__thisSynchronized    ;
  input                                         pe13__sys__ready               ;
  input                                         pe13__sys__complete            ;

  // General control and status                                                   
  input                                         mgr14__sys__allSynchronized     ;
  output                                        sys__mgr14__thisSynchronized    ;
  output                                        sys__mgr14__ready               ;
  output                                        sys__mgr14__complete            ;

  output                                        sys__pe14__allSynchronized     ;
  input                                         pe14__sys__thisSynchronized    ;
  input                                         pe14__sys__ready               ;
  input                                         pe14__sys__complete            ;

  // General control and status                                                   
  input                                         mgr15__sys__allSynchronized     ;
  output                                        sys__mgr15__thisSynchronized    ;
  output                                        sys__mgr15__ready               ;
  output                                        sys__mgr15__complete            ;

  output                                        sys__pe15__allSynchronized     ;
  input                                         pe15__sys__thisSynchronized    ;
  input                                         pe15__sys__ready               ;
  input                                         pe15__sys__complete            ;

  // General control and status                                                   
  input                                         mgr16__sys__allSynchronized     ;
  output                                        sys__mgr16__thisSynchronized    ;
  output                                        sys__mgr16__ready               ;
  output                                        sys__mgr16__complete            ;

  output                                        sys__pe16__allSynchronized     ;
  input                                         pe16__sys__thisSynchronized    ;
  input                                         pe16__sys__ready               ;
  input                                         pe16__sys__complete            ;

  // General control and status                                                   
  input                                         mgr17__sys__allSynchronized     ;
  output                                        sys__mgr17__thisSynchronized    ;
  output                                        sys__mgr17__ready               ;
  output                                        sys__mgr17__complete            ;

  output                                        sys__pe17__allSynchronized     ;
  input                                         pe17__sys__thisSynchronized    ;
  input                                         pe17__sys__ready               ;
  input                                         pe17__sys__complete            ;

  // General control and status                                                   
  input                                         mgr18__sys__allSynchronized     ;
  output                                        sys__mgr18__thisSynchronized    ;
  output                                        sys__mgr18__ready               ;
  output                                        sys__mgr18__complete            ;

  output                                        sys__pe18__allSynchronized     ;
  input                                         pe18__sys__thisSynchronized    ;
  input                                         pe18__sys__ready               ;
  input                                         pe18__sys__complete            ;

  // General control and status                                                   
  input                                         mgr19__sys__allSynchronized     ;
  output                                        sys__mgr19__thisSynchronized    ;
  output                                        sys__mgr19__ready               ;
  output                                        sys__mgr19__complete            ;

  output                                        sys__pe19__allSynchronized     ;
  input                                         pe19__sys__thisSynchronized    ;
  input                                         pe19__sys__ready               ;
  input                                         pe19__sys__complete            ;

  // General control and status                                                   
  input                                         mgr20__sys__allSynchronized     ;
  output                                        sys__mgr20__thisSynchronized    ;
  output                                        sys__mgr20__ready               ;
  output                                        sys__mgr20__complete            ;

  output                                        sys__pe20__allSynchronized     ;
  input                                         pe20__sys__thisSynchronized    ;
  input                                         pe20__sys__ready               ;
  input                                         pe20__sys__complete            ;

  // General control and status                                                   
  input                                         mgr21__sys__allSynchronized     ;
  output                                        sys__mgr21__thisSynchronized    ;
  output                                        sys__mgr21__ready               ;
  output                                        sys__mgr21__complete            ;

  output                                        sys__pe21__allSynchronized     ;
  input                                         pe21__sys__thisSynchronized    ;
  input                                         pe21__sys__ready               ;
  input                                         pe21__sys__complete            ;

  // General control and status                                                   
  input                                         mgr22__sys__allSynchronized     ;
  output                                        sys__mgr22__thisSynchronized    ;
  output                                        sys__mgr22__ready               ;
  output                                        sys__mgr22__complete            ;

  output                                        sys__pe22__allSynchronized     ;
  input                                         pe22__sys__thisSynchronized    ;
  input                                         pe22__sys__ready               ;
  input                                         pe22__sys__complete            ;

  // General control and status                                                   
  input                                         mgr23__sys__allSynchronized     ;
  output                                        sys__mgr23__thisSynchronized    ;
  output                                        sys__mgr23__ready               ;
  output                                        sys__mgr23__complete            ;

  output                                        sys__pe23__allSynchronized     ;
  input                                         pe23__sys__thisSynchronized    ;
  input                                         pe23__sys__ready               ;
  input                                         pe23__sys__complete            ;

  // General control and status                                                   
  input                                         mgr24__sys__allSynchronized     ;
  output                                        sys__mgr24__thisSynchronized    ;
  output                                        sys__mgr24__ready               ;
  output                                        sys__mgr24__complete            ;

  output                                        sys__pe24__allSynchronized     ;
  input                                         pe24__sys__thisSynchronized    ;
  input                                         pe24__sys__ready               ;
  input                                         pe24__sys__complete            ;

  // General control and status                                                   
  input                                         mgr25__sys__allSynchronized     ;
  output                                        sys__mgr25__thisSynchronized    ;
  output                                        sys__mgr25__ready               ;
  output                                        sys__mgr25__complete            ;

  output                                        sys__pe25__allSynchronized     ;
  input                                         pe25__sys__thisSynchronized    ;
  input                                         pe25__sys__ready               ;
  input                                         pe25__sys__complete            ;

  // General control and status                                                   
  input                                         mgr26__sys__allSynchronized     ;
  output                                        sys__mgr26__thisSynchronized    ;
  output                                        sys__mgr26__ready               ;
  output                                        sys__mgr26__complete            ;

  output                                        sys__pe26__allSynchronized     ;
  input                                         pe26__sys__thisSynchronized    ;
  input                                         pe26__sys__ready               ;
  input                                         pe26__sys__complete            ;

  // General control and status                                                   
  input                                         mgr27__sys__allSynchronized     ;
  output                                        sys__mgr27__thisSynchronized    ;
  output                                        sys__mgr27__ready               ;
  output                                        sys__mgr27__complete            ;

  output                                        sys__pe27__allSynchronized     ;
  input                                         pe27__sys__thisSynchronized    ;
  input                                         pe27__sys__ready               ;
  input                                         pe27__sys__complete            ;

  // General control and status                                                   
  input                                         mgr28__sys__allSynchronized     ;
  output                                        sys__mgr28__thisSynchronized    ;
  output                                        sys__mgr28__ready               ;
  output                                        sys__mgr28__complete            ;

  output                                        sys__pe28__allSynchronized     ;
  input                                         pe28__sys__thisSynchronized    ;
  input                                         pe28__sys__ready               ;
  input                                         pe28__sys__complete            ;

  // General control and status                                                   
  input                                         mgr29__sys__allSynchronized     ;
  output                                        sys__mgr29__thisSynchronized    ;
  output                                        sys__mgr29__ready               ;
  output                                        sys__mgr29__complete            ;

  output                                        sys__pe29__allSynchronized     ;
  input                                         pe29__sys__thisSynchronized    ;
  input                                         pe29__sys__ready               ;
  input                                         pe29__sys__complete            ;

  // General control and status                                                   
  input                                         mgr30__sys__allSynchronized     ;
  output                                        sys__mgr30__thisSynchronized    ;
  output                                        sys__mgr30__ready               ;
  output                                        sys__mgr30__complete            ;

  output                                        sys__pe30__allSynchronized     ;
  input                                         pe30__sys__thisSynchronized    ;
  input                                         pe30__sys__ready               ;
  input                                         pe30__sys__complete            ;

  // General control and status                                                   
  input                                         mgr31__sys__allSynchronized     ;
  output                                        sys__mgr31__thisSynchronized    ;
  output                                        sys__mgr31__ready               ;
  output                                        sys__mgr31__complete            ;

  output                                        sys__pe31__allSynchronized     ;
  input                                         pe31__sys__thisSynchronized    ;
  input                                         pe31__sys__ready               ;
  input                                         pe31__sys__complete            ;

  // General control and status                                                   
  input                                         mgr32__sys__allSynchronized     ;
  output                                        sys__mgr32__thisSynchronized    ;
  output                                        sys__mgr32__ready               ;
  output                                        sys__mgr32__complete            ;

  output                                        sys__pe32__allSynchronized     ;
  input                                         pe32__sys__thisSynchronized    ;
  input                                         pe32__sys__ready               ;
  input                                         pe32__sys__complete            ;

  // General control and status                                                   
  input                                         mgr33__sys__allSynchronized     ;
  output                                        sys__mgr33__thisSynchronized    ;
  output                                        sys__mgr33__ready               ;
  output                                        sys__mgr33__complete            ;

  output                                        sys__pe33__allSynchronized     ;
  input                                         pe33__sys__thisSynchronized    ;
  input                                         pe33__sys__ready               ;
  input                                         pe33__sys__complete            ;

  // General control and status                                                   
  input                                         mgr34__sys__allSynchronized     ;
  output                                        sys__mgr34__thisSynchronized    ;
  output                                        sys__mgr34__ready               ;
  output                                        sys__mgr34__complete            ;

  output                                        sys__pe34__allSynchronized     ;
  input                                         pe34__sys__thisSynchronized    ;
  input                                         pe34__sys__ready               ;
  input                                         pe34__sys__complete            ;

  // General control and status                                                   
  input                                         mgr35__sys__allSynchronized     ;
  output                                        sys__mgr35__thisSynchronized    ;
  output                                        sys__mgr35__ready               ;
  output                                        sys__mgr35__complete            ;

  output                                        sys__pe35__allSynchronized     ;
  input                                         pe35__sys__thisSynchronized    ;
  input                                         pe35__sys__ready               ;
  input                                         pe35__sys__complete            ;

  // General control and status                                                   
  input                                         mgr36__sys__allSynchronized     ;
  output                                        sys__mgr36__thisSynchronized    ;
  output                                        sys__mgr36__ready               ;
  output                                        sys__mgr36__complete            ;

  output                                        sys__pe36__allSynchronized     ;
  input                                         pe36__sys__thisSynchronized    ;
  input                                         pe36__sys__ready               ;
  input                                         pe36__sys__complete            ;

  // General control and status                                                   
  input                                         mgr37__sys__allSynchronized     ;
  output                                        sys__mgr37__thisSynchronized    ;
  output                                        sys__mgr37__ready               ;
  output                                        sys__mgr37__complete            ;

  output                                        sys__pe37__allSynchronized     ;
  input                                         pe37__sys__thisSynchronized    ;
  input                                         pe37__sys__ready               ;
  input                                         pe37__sys__complete            ;

  // General control and status                                                   
  input                                         mgr38__sys__allSynchronized     ;
  output                                        sys__mgr38__thisSynchronized    ;
  output                                        sys__mgr38__ready               ;
  output                                        sys__mgr38__complete            ;

  output                                        sys__pe38__allSynchronized     ;
  input                                         pe38__sys__thisSynchronized    ;
  input                                         pe38__sys__ready               ;
  input                                         pe38__sys__complete            ;

  // General control and status                                                   
  input                                         mgr39__sys__allSynchronized     ;
  output                                        sys__mgr39__thisSynchronized    ;
  output                                        sys__mgr39__ready               ;
  output                                        sys__mgr39__complete            ;

  output                                        sys__pe39__allSynchronized     ;
  input                                         pe39__sys__thisSynchronized    ;
  input                                         pe39__sys__ready               ;
  input                                         pe39__sys__complete            ;

  // General control and status                                                   
  input                                         mgr40__sys__allSynchronized     ;
  output                                        sys__mgr40__thisSynchronized    ;
  output                                        sys__mgr40__ready               ;
  output                                        sys__mgr40__complete            ;

  output                                        sys__pe40__allSynchronized     ;
  input                                         pe40__sys__thisSynchronized    ;
  input                                         pe40__sys__ready               ;
  input                                         pe40__sys__complete            ;

  // General control and status                                                   
  input                                         mgr41__sys__allSynchronized     ;
  output                                        sys__mgr41__thisSynchronized    ;
  output                                        sys__mgr41__ready               ;
  output                                        sys__mgr41__complete            ;

  output                                        sys__pe41__allSynchronized     ;
  input                                         pe41__sys__thisSynchronized    ;
  input                                         pe41__sys__ready               ;
  input                                         pe41__sys__complete            ;

  // General control and status                                                   
  input                                         mgr42__sys__allSynchronized     ;
  output                                        sys__mgr42__thisSynchronized    ;
  output                                        sys__mgr42__ready               ;
  output                                        sys__mgr42__complete            ;

  output                                        sys__pe42__allSynchronized     ;
  input                                         pe42__sys__thisSynchronized    ;
  input                                         pe42__sys__ready               ;
  input                                         pe42__sys__complete            ;

  // General control and status                                                   
  input                                         mgr43__sys__allSynchronized     ;
  output                                        sys__mgr43__thisSynchronized    ;
  output                                        sys__mgr43__ready               ;
  output                                        sys__mgr43__complete            ;

  output                                        sys__pe43__allSynchronized     ;
  input                                         pe43__sys__thisSynchronized    ;
  input                                         pe43__sys__ready               ;
  input                                         pe43__sys__complete            ;

  // General control and status                                                   
  input                                         mgr44__sys__allSynchronized     ;
  output                                        sys__mgr44__thisSynchronized    ;
  output                                        sys__mgr44__ready               ;
  output                                        sys__mgr44__complete            ;

  output                                        sys__pe44__allSynchronized     ;
  input                                         pe44__sys__thisSynchronized    ;
  input                                         pe44__sys__ready               ;
  input                                         pe44__sys__complete            ;

  // General control and status                                                   
  input                                         mgr45__sys__allSynchronized     ;
  output                                        sys__mgr45__thisSynchronized    ;
  output                                        sys__mgr45__ready               ;
  output                                        sys__mgr45__complete            ;

  output                                        sys__pe45__allSynchronized     ;
  input                                         pe45__sys__thisSynchronized    ;
  input                                         pe45__sys__ready               ;
  input                                         pe45__sys__complete            ;

  // General control and status                                                   
  input                                         mgr46__sys__allSynchronized     ;
  output                                        sys__mgr46__thisSynchronized    ;
  output                                        sys__mgr46__ready               ;
  output                                        sys__mgr46__complete            ;

  output                                        sys__pe46__allSynchronized     ;
  input                                         pe46__sys__thisSynchronized    ;
  input                                         pe46__sys__ready               ;
  input                                         pe46__sys__complete            ;

  // General control and status                                                   
  input                                         mgr47__sys__allSynchronized     ;
  output                                        sys__mgr47__thisSynchronized    ;
  output                                        sys__mgr47__ready               ;
  output                                        sys__mgr47__complete            ;

  output                                        sys__pe47__allSynchronized     ;
  input                                         pe47__sys__thisSynchronized    ;
  input                                         pe47__sys__ready               ;
  input                                         pe47__sys__complete            ;

  // General control and status                                                   
  input                                         mgr48__sys__allSynchronized     ;
  output                                        sys__mgr48__thisSynchronized    ;
  output                                        sys__mgr48__ready               ;
  output                                        sys__mgr48__complete            ;

  output                                        sys__pe48__allSynchronized     ;
  input                                         pe48__sys__thisSynchronized    ;
  input                                         pe48__sys__ready               ;
  input                                         pe48__sys__complete            ;

  // General control and status                                                   
  input                                         mgr49__sys__allSynchronized     ;
  output                                        sys__mgr49__thisSynchronized    ;
  output                                        sys__mgr49__ready               ;
  output                                        sys__mgr49__complete            ;

  output                                        sys__pe49__allSynchronized     ;
  input                                         pe49__sys__thisSynchronized    ;
  input                                         pe49__sys__ready               ;
  input                                         pe49__sys__complete            ;

  // General control and status                                                   
  input                                         mgr50__sys__allSynchronized     ;
  output                                        sys__mgr50__thisSynchronized    ;
  output                                        sys__mgr50__ready               ;
  output                                        sys__mgr50__complete            ;

  output                                        sys__pe50__allSynchronized     ;
  input                                         pe50__sys__thisSynchronized    ;
  input                                         pe50__sys__ready               ;
  input                                         pe50__sys__complete            ;

  // General control and status                                                   
  input                                         mgr51__sys__allSynchronized     ;
  output                                        sys__mgr51__thisSynchronized    ;
  output                                        sys__mgr51__ready               ;
  output                                        sys__mgr51__complete            ;

  output                                        sys__pe51__allSynchronized     ;
  input                                         pe51__sys__thisSynchronized    ;
  input                                         pe51__sys__ready               ;
  input                                         pe51__sys__complete            ;

  // General control and status                                                   
  input                                         mgr52__sys__allSynchronized     ;
  output                                        sys__mgr52__thisSynchronized    ;
  output                                        sys__mgr52__ready               ;
  output                                        sys__mgr52__complete            ;

  output                                        sys__pe52__allSynchronized     ;
  input                                         pe52__sys__thisSynchronized    ;
  input                                         pe52__sys__ready               ;
  input                                         pe52__sys__complete            ;

  // General control and status                                                   
  input                                         mgr53__sys__allSynchronized     ;
  output                                        sys__mgr53__thisSynchronized    ;
  output                                        sys__mgr53__ready               ;
  output                                        sys__mgr53__complete            ;

  output                                        sys__pe53__allSynchronized     ;
  input                                         pe53__sys__thisSynchronized    ;
  input                                         pe53__sys__ready               ;
  input                                         pe53__sys__complete            ;

  // General control and status                                                   
  input                                         mgr54__sys__allSynchronized     ;
  output                                        sys__mgr54__thisSynchronized    ;
  output                                        sys__mgr54__ready               ;
  output                                        sys__mgr54__complete            ;

  output                                        sys__pe54__allSynchronized     ;
  input                                         pe54__sys__thisSynchronized    ;
  input                                         pe54__sys__ready               ;
  input                                         pe54__sys__complete            ;

  // General control and status                                                   
  input                                         mgr55__sys__allSynchronized     ;
  output                                        sys__mgr55__thisSynchronized    ;
  output                                        sys__mgr55__ready               ;
  output                                        sys__mgr55__complete            ;

  output                                        sys__pe55__allSynchronized     ;
  input                                         pe55__sys__thisSynchronized    ;
  input                                         pe55__sys__ready               ;
  input                                         pe55__sys__complete            ;

  // General control and status                                                   
  input                                         mgr56__sys__allSynchronized     ;
  output                                        sys__mgr56__thisSynchronized    ;
  output                                        sys__mgr56__ready               ;
  output                                        sys__mgr56__complete            ;

  output                                        sys__pe56__allSynchronized     ;
  input                                         pe56__sys__thisSynchronized    ;
  input                                         pe56__sys__ready               ;
  input                                         pe56__sys__complete            ;

  // General control and status                                                   
  input                                         mgr57__sys__allSynchronized     ;
  output                                        sys__mgr57__thisSynchronized    ;
  output                                        sys__mgr57__ready               ;
  output                                        sys__mgr57__complete            ;

  output                                        sys__pe57__allSynchronized     ;
  input                                         pe57__sys__thisSynchronized    ;
  input                                         pe57__sys__ready               ;
  input                                         pe57__sys__complete            ;

  // General control and status                                                   
  input                                         mgr58__sys__allSynchronized     ;
  output                                        sys__mgr58__thisSynchronized    ;
  output                                        sys__mgr58__ready               ;
  output                                        sys__mgr58__complete            ;

  output                                        sys__pe58__allSynchronized     ;
  input                                         pe58__sys__thisSynchronized    ;
  input                                         pe58__sys__ready               ;
  input                                         pe58__sys__complete            ;

  // General control and status                                                   
  input                                         mgr59__sys__allSynchronized     ;
  output                                        sys__mgr59__thisSynchronized    ;
  output                                        sys__mgr59__ready               ;
  output                                        sys__mgr59__complete            ;

  output                                        sys__pe59__allSynchronized     ;
  input                                         pe59__sys__thisSynchronized    ;
  input                                         pe59__sys__ready               ;
  input                                         pe59__sys__complete            ;

  // General control and status                                                   
  input                                         mgr60__sys__allSynchronized     ;
  output                                        sys__mgr60__thisSynchronized    ;
  output                                        sys__mgr60__ready               ;
  output                                        sys__mgr60__complete            ;

  output                                        sys__pe60__allSynchronized     ;
  input                                         pe60__sys__thisSynchronized    ;
  input                                         pe60__sys__ready               ;
  input                                         pe60__sys__complete            ;

  // General control and status                                                   
  input                                         mgr61__sys__allSynchronized     ;
  output                                        sys__mgr61__thisSynchronized    ;
  output                                        sys__mgr61__ready               ;
  output                                        sys__mgr61__complete            ;

  output                                        sys__pe61__allSynchronized     ;
  input                                         pe61__sys__thisSynchronized    ;
  input                                         pe61__sys__ready               ;
  input                                         pe61__sys__complete            ;

  // General control and status                                                   
  input                                         mgr62__sys__allSynchronized     ;
  output                                        sys__mgr62__thisSynchronized    ;
  output                                        sys__mgr62__ready               ;
  output                                        sys__mgr62__complete            ;

  output                                        sys__pe62__allSynchronized     ;
  input                                         pe62__sys__thisSynchronized    ;
  input                                         pe62__sys__ready               ;
  input                                         pe62__sys__complete            ;

  // General control and status                                                   
  input                                         mgr63__sys__allSynchronized     ;
  output                                        sys__mgr63__thisSynchronized    ;
  output                                        sys__mgr63__ready               ;
  output                                        sys__mgr63__complete            ;

  output                                        sys__pe63__allSynchronized     ;
  input                                         pe63__sys__thisSynchronized    ;
  input                                         pe63__sys__ready               ;
  input                                         pe63__sys__complete            ;
