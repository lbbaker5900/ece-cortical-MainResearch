
  output                                    reg__scntl__lane0_ready    ;
  input                                     scntl__reg__lane0_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane0_data     ;

  output                                    reg__scntl__lane1_ready    ;
  input                                     scntl__reg__lane1_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane1_data     ;

  output                                    reg__scntl__lane2_ready    ;
  input                                     scntl__reg__lane2_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane2_data     ;

  output                                    reg__scntl__lane3_ready    ;
  input                                     scntl__reg__lane3_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane3_data     ;

  output                                    reg__scntl__lane4_ready    ;
  input                                     scntl__reg__lane4_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane4_data     ;

  output                                    reg__scntl__lane5_ready    ;
  input                                     scntl__reg__lane5_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane5_data     ;

  output                                    reg__scntl__lane6_ready    ;
  input                                     scntl__reg__lane6_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane6_data     ;

  output                                    reg__scntl__lane7_ready    ;
  input                                     scntl__reg__lane7_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane7_data     ;

  output                                    reg__scntl__lane8_ready    ;
  input                                     scntl__reg__lane8_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane8_data     ;

  output                                    reg__scntl__lane9_ready    ;
  input                                     scntl__reg__lane9_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane9_data     ;

  output                                    reg__scntl__lane10_ready    ;
  input                                     scntl__reg__lane10_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane10_data     ;

  output                                    reg__scntl__lane11_ready    ;
  input                                     scntl__reg__lane11_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane11_data     ;

  output                                    reg__scntl__lane12_ready    ;
  input                                     scntl__reg__lane12_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane12_data     ;

  output                                    reg__scntl__lane13_ready    ;
  input                                     scntl__reg__lane13_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane13_data     ;

  output                                    reg__scntl__lane14_ready    ;
  input                                     scntl__reg__lane14_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane14_data     ;

  output                                    reg__scntl__lane15_ready    ;
  input                                     scntl__reg__lane15_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane15_data     ;

  output                                    reg__scntl__lane16_ready    ;
  input                                     scntl__reg__lane16_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane16_data     ;

  output                                    reg__scntl__lane17_ready    ;
  input                                     scntl__reg__lane17_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane17_data     ;

  output                                    reg__scntl__lane18_ready    ;
  input                                     scntl__reg__lane18_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane18_data     ;

  output                                    reg__scntl__lane19_ready    ;
  input                                     scntl__reg__lane19_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane19_data     ;

  output                                    reg__scntl__lane20_ready    ;
  input                                     scntl__reg__lane20_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane20_data     ;

  output                                    reg__scntl__lane21_ready    ;
  input                                     scntl__reg__lane21_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane21_data     ;

  output                                    reg__scntl__lane22_ready    ;
  input                                     scntl__reg__lane22_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane22_data     ;

  output                                    reg__scntl__lane23_ready    ;
  input                                     scntl__reg__lane23_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane23_data     ;

  output                                    reg__scntl__lane24_ready    ;
  input                                     scntl__reg__lane24_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane24_data     ;

  output                                    reg__scntl__lane25_ready    ;
  input                                     scntl__reg__lane25_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane25_data     ;

  output                                    reg__scntl__lane26_ready    ;
  input                                     scntl__reg__lane26_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane26_data     ;

  output                                    reg__scntl__lane27_ready    ;
  input                                     scntl__reg__lane27_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane27_data     ;

  output                                    reg__scntl__lane28_ready    ;
  input                                     scntl__reg__lane28_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane28_data     ;

  output                                    reg__scntl__lane29_ready    ;
  input                                     scntl__reg__lane29_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane29_data     ;

  output                                    reg__scntl__lane30_ready    ;
  input                                     scntl__reg__lane30_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane30_data     ;

  output                                    reg__scntl__lane31_ready    ;
  input                                     scntl__reg__lane31_valid    ;
  input    [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane31_data     ;

