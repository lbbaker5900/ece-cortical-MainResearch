
            begin
              mr_proc[0][0].run()  ;
            end

            begin
              mr_proc[0][1].run()  ;
            end

            begin
              mr_proc[1][0].run()  ;
            end

            begin
              mr_proc[1][1].run()  ;
            end

            begin
              mr_proc[2][0].run()  ;
            end

            begin
              mr_proc[2][1].run()  ;
            end

            begin
              mr_proc[3][0].run()  ;
            end

            begin
              mr_proc[3][1].run()  ;
            end
