
            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 0, lane 0, stream 0      
            input   wire                                        std__mgr0__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane0_strm0_data        ,
            output  wire                                        mgr0__std__lane0_strm0_data_valid  ,

            // manager 0, lane 0, stream 1      
            input   wire                                        std__mgr0__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane0_strm1_data        ,
            output  wire                                        mgr0__std__lane0_strm1_data_valid  ,

            // manager 0, lane 1, stream 0      
            input   wire                                        std__mgr0__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane1_strm0_data        ,
            output  wire                                        mgr0__std__lane1_strm0_data_valid  ,

            // manager 0, lane 1, stream 1      
            input   wire                                        std__mgr0__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane1_strm1_data        ,
            output  wire                                        mgr0__std__lane1_strm1_data_valid  ,

            // manager 0, lane 2, stream 0      
            input   wire                                        std__mgr0__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane2_strm0_data        ,
            output  wire                                        mgr0__std__lane2_strm0_data_valid  ,

            // manager 0, lane 2, stream 1      
            input   wire                                        std__mgr0__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane2_strm1_data        ,
            output  wire                                        mgr0__std__lane2_strm1_data_valid  ,

            // manager 0, lane 3, stream 0      
            input   wire                                        std__mgr0__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane3_strm0_data        ,
            output  wire                                        mgr0__std__lane3_strm0_data_valid  ,

            // manager 0, lane 3, stream 1      
            input   wire                                        std__mgr0__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane3_strm1_data        ,
            output  wire                                        mgr0__std__lane3_strm1_data_valid  ,

            // manager 0, lane 4, stream 0      
            input   wire                                        std__mgr0__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane4_strm0_data        ,
            output  wire                                        mgr0__std__lane4_strm0_data_valid  ,

            // manager 0, lane 4, stream 1      
            input   wire                                        std__mgr0__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane4_strm1_data        ,
            output  wire                                        mgr0__std__lane4_strm1_data_valid  ,

            // manager 0, lane 5, stream 0      
            input   wire                                        std__mgr0__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane5_strm0_data        ,
            output  wire                                        mgr0__std__lane5_strm0_data_valid  ,

            // manager 0, lane 5, stream 1      
            input   wire                                        std__mgr0__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane5_strm1_data        ,
            output  wire                                        mgr0__std__lane5_strm1_data_valid  ,

            // manager 0, lane 6, stream 0      
            input   wire                                        std__mgr0__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane6_strm0_data        ,
            output  wire                                        mgr0__std__lane6_strm0_data_valid  ,

            // manager 0, lane 6, stream 1      
            input   wire                                        std__mgr0__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane6_strm1_data        ,
            output  wire                                        mgr0__std__lane6_strm1_data_valid  ,

            // manager 0, lane 7, stream 0      
            input   wire                                        std__mgr0__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane7_strm0_data        ,
            output  wire                                        mgr0__std__lane7_strm0_data_valid  ,

            // manager 0, lane 7, stream 1      
            input   wire                                        std__mgr0__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane7_strm1_data        ,
            output  wire                                        mgr0__std__lane7_strm1_data_valid  ,

            // manager 0, lane 8, stream 0      
            input   wire                                        std__mgr0__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane8_strm0_data        ,
            output  wire                                        mgr0__std__lane8_strm0_data_valid  ,

            // manager 0, lane 8, stream 1      
            input   wire                                        std__mgr0__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane8_strm1_data        ,
            output  wire                                        mgr0__std__lane8_strm1_data_valid  ,

            // manager 0, lane 9, stream 0      
            input   wire                                        std__mgr0__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane9_strm0_data        ,
            output  wire                                        mgr0__std__lane9_strm0_data_valid  ,

            // manager 0, lane 9, stream 1      
            input   wire                                        std__mgr0__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane9_strm1_data        ,
            output  wire                                        mgr0__std__lane9_strm1_data_valid  ,

            // manager 0, lane 10, stream 0      
            input   wire                                        std__mgr0__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane10_strm0_data        ,
            output  wire                                        mgr0__std__lane10_strm0_data_valid  ,

            // manager 0, lane 10, stream 1      
            input   wire                                        std__mgr0__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane10_strm1_data        ,
            output  wire                                        mgr0__std__lane10_strm1_data_valid  ,

            // manager 0, lane 11, stream 0      
            input   wire                                        std__mgr0__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane11_strm0_data        ,
            output  wire                                        mgr0__std__lane11_strm0_data_valid  ,

            // manager 0, lane 11, stream 1      
            input   wire                                        std__mgr0__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane11_strm1_data        ,
            output  wire                                        mgr0__std__lane11_strm1_data_valid  ,

            // manager 0, lane 12, stream 0      
            input   wire                                        std__mgr0__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane12_strm0_data        ,
            output  wire                                        mgr0__std__lane12_strm0_data_valid  ,

            // manager 0, lane 12, stream 1      
            input   wire                                        std__mgr0__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane12_strm1_data        ,
            output  wire                                        mgr0__std__lane12_strm1_data_valid  ,

            // manager 0, lane 13, stream 0      
            input   wire                                        std__mgr0__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane13_strm0_data        ,
            output  wire                                        mgr0__std__lane13_strm0_data_valid  ,

            // manager 0, lane 13, stream 1      
            input   wire                                        std__mgr0__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane13_strm1_data        ,
            output  wire                                        mgr0__std__lane13_strm1_data_valid  ,

            // manager 0, lane 14, stream 0      
            input   wire                                        std__mgr0__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane14_strm0_data        ,
            output  wire                                        mgr0__std__lane14_strm0_data_valid  ,

            // manager 0, lane 14, stream 1      
            input   wire                                        std__mgr0__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane14_strm1_data        ,
            output  wire                                        mgr0__std__lane14_strm1_data_valid  ,

            // manager 0, lane 15, stream 0      
            input   wire                                        std__mgr0__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane15_strm0_data        ,
            output  wire                                        mgr0__std__lane15_strm0_data_valid  ,

            // manager 0, lane 15, stream 1      
            input   wire                                        std__mgr0__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane15_strm1_data        ,
            output  wire                                        mgr0__std__lane15_strm1_data_valid  ,

            // manager 0, lane 16, stream 0      
            input   wire                                        std__mgr0__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane16_strm0_data        ,
            output  wire                                        mgr0__std__lane16_strm0_data_valid  ,

            // manager 0, lane 16, stream 1      
            input   wire                                        std__mgr0__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane16_strm1_data        ,
            output  wire                                        mgr0__std__lane16_strm1_data_valid  ,

            // manager 0, lane 17, stream 0      
            input   wire                                        std__mgr0__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane17_strm0_data        ,
            output  wire                                        mgr0__std__lane17_strm0_data_valid  ,

            // manager 0, lane 17, stream 1      
            input   wire                                        std__mgr0__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane17_strm1_data        ,
            output  wire                                        mgr0__std__lane17_strm1_data_valid  ,

            // manager 0, lane 18, stream 0      
            input   wire                                        std__mgr0__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane18_strm0_data        ,
            output  wire                                        mgr0__std__lane18_strm0_data_valid  ,

            // manager 0, lane 18, stream 1      
            input   wire                                        std__mgr0__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane18_strm1_data        ,
            output  wire                                        mgr0__std__lane18_strm1_data_valid  ,

            // manager 0, lane 19, stream 0      
            input   wire                                        std__mgr0__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane19_strm0_data        ,
            output  wire                                        mgr0__std__lane19_strm0_data_valid  ,

            // manager 0, lane 19, stream 1      
            input   wire                                        std__mgr0__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane19_strm1_data        ,
            output  wire                                        mgr0__std__lane19_strm1_data_valid  ,

            // manager 0, lane 20, stream 0      
            input   wire                                        std__mgr0__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane20_strm0_data        ,
            output  wire                                        mgr0__std__lane20_strm0_data_valid  ,

            // manager 0, lane 20, stream 1      
            input   wire                                        std__mgr0__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane20_strm1_data        ,
            output  wire                                        mgr0__std__lane20_strm1_data_valid  ,

            // manager 0, lane 21, stream 0      
            input   wire                                        std__mgr0__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane21_strm0_data        ,
            output  wire                                        mgr0__std__lane21_strm0_data_valid  ,

            // manager 0, lane 21, stream 1      
            input   wire                                        std__mgr0__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane21_strm1_data        ,
            output  wire                                        mgr0__std__lane21_strm1_data_valid  ,

            // manager 0, lane 22, stream 0      
            input   wire                                        std__mgr0__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane22_strm0_data        ,
            output  wire                                        mgr0__std__lane22_strm0_data_valid  ,

            // manager 0, lane 22, stream 1      
            input   wire                                        std__mgr0__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane22_strm1_data        ,
            output  wire                                        mgr0__std__lane22_strm1_data_valid  ,

            // manager 0, lane 23, stream 0      
            input   wire                                        std__mgr0__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane23_strm0_data        ,
            output  wire                                        mgr0__std__lane23_strm0_data_valid  ,

            // manager 0, lane 23, stream 1      
            input   wire                                        std__mgr0__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane23_strm1_data        ,
            output  wire                                        mgr0__std__lane23_strm1_data_valid  ,

            // manager 0, lane 24, stream 0      
            input   wire                                        std__mgr0__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane24_strm0_data        ,
            output  wire                                        mgr0__std__lane24_strm0_data_valid  ,

            // manager 0, lane 24, stream 1      
            input   wire                                        std__mgr0__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane24_strm1_data        ,
            output  wire                                        mgr0__std__lane24_strm1_data_valid  ,

            // manager 0, lane 25, stream 0      
            input   wire                                        std__mgr0__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane25_strm0_data        ,
            output  wire                                        mgr0__std__lane25_strm0_data_valid  ,

            // manager 0, lane 25, stream 1      
            input   wire                                        std__mgr0__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane25_strm1_data        ,
            output  wire                                        mgr0__std__lane25_strm1_data_valid  ,

            // manager 0, lane 26, stream 0      
            input   wire                                        std__mgr0__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane26_strm0_data        ,
            output  wire                                        mgr0__std__lane26_strm0_data_valid  ,

            // manager 0, lane 26, stream 1      
            input   wire                                        std__mgr0__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane26_strm1_data        ,
            output  wire                                        mgr0__std__lane26_strm1_data_valid  ,

            // manager 0, lane 27, stream 0      
            input   wire                                        std__mgr0__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane27_strm0_data        ,
            output  wire                                        mgr0__std__lane27_strm0_data_valid  ,

            // manager 0, lane 27, stream 1      
            input   wire                                        std__mgr0__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane27_strm1_data        ,
            output  wire                                        mgr0__std__lane27_strm1_data_valid  ,

            // manager 0, lane 28, stream 0      
            input   wire                                        std__mgr0__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane28_strm0_data        ,
            output  wire                                        mgr0__std__lane28_strm0_data_valid  ,

            // manager 0, lane 28, stream 1      
            input   wire                                        std__mgr0__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane28_strm1_data        ,
            output  wire                                        mgr0__std__lane28_strm1_data_valid  ,

            // manager 0, lane 29, stream 0      
            input   wire                                        std__mgr0__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane29_strm0_data        ,
            output  wire                                        mgr0__std__lane29_strm0_data_valid  ,

            // manager 0, lane 29, stream 1      
            input   wire                                        std__mgr0__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane29_strm1_data        ,
            output  wire                                        mgr0__std__lane29_strm1_data_valid  ,

            // manager 0, lane 30, stream 0      
            input   wire                                        std__mgr0__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane30_strm0_data        ,
            output  wire                                        mgr0__std__lane30_strm0_data_valid  ,

            // manager 0, lane 30, stream 1      
            input   wire                                        std__mgr0__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane30_strm1_data        ,
            output  wire                                        mgr0__std__lane30_strm1_data_valid  ,

            // manager 0, lane 31, stream 0      
            input   wire                                        std__mgr0__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane31_strm0_data        ,
            output  wire                                        mgr0__std__lane31_strm0_data_valid  ,

            // manager 0, lane 31, stream 1      
            input   wire                                        std__mgr0__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr0__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr0__std__lane31_strm1_data        ,
            output  wire                                        mgr0__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 1, lane 0, stream 0      
            input   wire                                        std__mgr1__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane0_strm0_data        ,
            output  wire                                        mgr1__std__lane0_strm0_data_valid  ,

            // manager 1, lane 0, stream 1      
            input   wire                                        std__mgr1__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane0_strm1_data        ,
            output  wire                                        mgr1__std__lane0_strm1_data_valid  ,

            // manager 1, lane 1, stream 0      
            input   wire                                        std__mgr1__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane1_strm0_data        ,
            output  wire                                        mgr1__std__lane1_strm0_data_valid  ,

            // manager 1, lane 1, stream 1      
            input   wire                                        std__mgr1__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane1_strm1_data        ,
            output  wire                                        mgr1__std__lane1_strm1_data_valid  ,

            // manager 1, lane 2, stream 0      
            input   wire                                        std__mgr1__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane2_strm0_data        ,
            output  wire                                        mgr1__std__lane2_strm0_data_valid  ,

            // manager 1, lane 2, stream 1      
            input   wire                                        std__mgr1__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane2_strm1_data        ,
            output  wire                                        mgr1__std__lane2_strm1_data_valid  ,

            // manager 1, lane 3, stream 0      
            input   wire                                        std__mgr1__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane3_strm0_data        ,
            output  wire                                        mgr1__std__lane3_strm0_data_valid  ,

            // manager 1, lane 3, stream 1      
            input   wire                                        std__mgr1__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane3_strm1_data        ,
            output  wire                                        mgr1__std__lane3_strm1_data_valid  ,

            // manager 1, lane 4, stream 0      
            input   wire                                        std__mgr1__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane4_strm0_data        ,
            output  wire                                        mgr1__std__lane4_strm0_data_valid  ,

            // manager 1, lane 4, stream 1      
            input   wire                                        std__mgr1__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane4_strm1_data        ,
            output  wire                                        mgr1__std__lane4_strm1_data_valid  ,

            // manager 1, lane 5, stream 0      
            input   wire                                        std__mgr1__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane5_strm0_data        ,
            output  wire                                        mgr1__std__lane5_strm0_data_valid  ,

            // manager 1, lane 5, stream 1      
            input   wire                                        std__mgr1__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane5_strm1_data        ,
            output  wire                                        mgr1__std__lane5_strm1_data_valid  ,

            // manager 1, lane 6, stream 0      
            input   wire                                        std__mgr1__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane6_strm0_data        ,
            output  wire                                        mgr1__std__lane6_strm0_data_valid  ,

            // manager 1, lane 6, stream 1      
            input   wire                                        std__mgr1__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane6_strm1_data        ,
            output  wire                                        mgr1__std__lane6_strm1_data_valid  ,

            // manager 1, lane 7, stream 0      
            input   wire                                        std__mgr1__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane7_strm0_data        ,
            output  wire                                        mgr1__std__lane7_strm0_data_valid  ,

            // manager 1, lane 7, stream 1      
            input   wire                                        std__mgr1__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane7_strm1_data        ,
            output  wire                                        mgr1__std__lane7_strm1_data_valid  ,

            // manager 1, lane 8, stream 0      
            input   wire                                        std__mgr1__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane8_strm0_data        ,
            output  wire                                        mgr1__std__lane8_strm0_data_valid  ,

            // manager 1, lane 8, stream 1      
            input   wire                                        std__mgr1__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane8_strm1_data        ,
            output  wire                                        mgr1__std__lane8_strm1_data_valid  ,

            // manager 1, lane 9, stream 0      
            input   wire                                        std__mgr1__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane9_strm0_data        ,
            output  wire                                        mgr1__std__lane9_strm0_data_valid  ,

            // manager 1, lane 9, stream 1      
            input   wire                                        std__mgr1__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane9_strm1_data        ,
            output  wire                                        mgr1__std__lane9_strm1_data_valid  ,

            // manager 1, lane 10, stream 0      
            input   wire                                        std__mgr1__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane10_strm0_data        ,
            output  wire                                        mgr1__std__lane10_strm0_data_valid  ,

            // manager 1, lane 10, stream 1      
            input   wire                                        std__mgr1__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane10_strm1_data        ,
            output  wire                                        mgr1__std__lane10_strm1_data_valid  ,

            // manager 1, lane 11, stream 0      
            input   wire                                        std__mgr1__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane11_strm0_data        ,
            output  wire                                        mgr1__std__lane11_strm0_data_valid  ,

            // manager 1, lane 11, stream 1      
            input   wire                                        std__mgr1__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane11_strm1_data        ,
            output  wire                                        mgr1__std__lane11_strm1_data_valid  ,

            // manager 1, lane 12, stream 0      
            input   wire                                        std__mgr1__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane12_strm0_data        ,
            output  wire                                        mgr1__std__lane12_strm0_data_valid  ,

            // manager 1, lane 12, stream 1      
            input   wire                                        std__mgr1__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane12_strm1_data        ,
            output  wire                                        mgr1__std__lane12_strm1_data_valid  ,

            // manager 1, lane 13, stream 0      
            input   wire                                        std__mgr1__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane13_strm0_data        ,
            output  wire                                        mgr1__std__lane13_strm0_data_valid  ,

            // manager 1, lane 13, stream 1      
            input   wire                                        std__mgr1__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane13_strm1_data        ,
            output  wire                                        mgr1__std__lane13_strm1_data_valid  ,

            // manager 1, lane 14, stream 0      
            input   wire                                        std__mgr1__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane14_strm0_data        ,
            output  wire                                        mgr1__std__lane14_strm0_data_valid  ,

            // manager 1, lane 14, stream 1      
            input   wire                                        std__mgr1__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane14_strm1_data        ,
            output  wire                                        mgr1__std__lane14_strm1_data_valid  ,

            // manager 1, lane 15, stream 0      
            input   wire                                        std__mgr1__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane15_strm0_data        ,
            output  wire                                        mgr1__std__lane15_strm0_data_valid  ,

            // manager 1, lane 15, stream 1      
            input   wire                                        std__mgr1__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane15_strm1_data        ,
            output  wire                                        mgr1__std__lane15_strm1_data_valid  ,

            // manager 1, lane 16, stream 0      
            input   wire                                        std__mgr1__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane16_strm0_data        ,
            output  wire                                        mgr1__std__lane16_strm0_data_valid  ,

            // manager 1, lane 16, stream 1      
            input   wire                                        std__mgr1__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane16_strm1_data        ,
            output  wire                                        mgr1__std__lane16_strm1_data_valid  ,

            // manager 1, lane 17, stream 0      
            input   wire                                        std__mgr1__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane17_strm0_data        ,
            output  wire                                        mgr1__std__lane17_strm0_data_valid  ,

            // manager 1, lane 17, stream 1      
            input   wire                                        std__mgr1__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane17_strm1_data        ,
            output  wire                                        mgr1__std__lane17_strm1_data_valid  ,

            // manager 1, lane 18, stream 0      
            input   wire                                        std__mgr1__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane18_strm0_data        ,
            output  wire                                        mgr1__std__lane18_strm0_data_valid  ,

            // manager 1, lane 18, stream 1      
            input   wire                                        std__mgr1__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane18_strm1_data        ,
            output  wire                                        mgr1__std__lane18_strm1_data_valid  ,

            // manager 1, lane 19, stream 0      
            input   wire                                        std__mgr1__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane19_strm0_data        ,
            output  wire                                        mgr1__std__lane19_strm0_data_valid  ,

            // manager 1, lane 19, stream 1      
            input   wire                                        std__mgr1__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane19_strm1_data        ,
            output  wire                                        mgr1__std__lane19_strm1_data_valid  ,

            // manager 1, lane 20, stream 0      
            input   wire                                        std__mgr1__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane20_strm0_data        ,
            output  wire                                        mgr1__std__lane20_strm0_data_valid  ,

            // manager 1, lane 20, stream 1      
            input   wire                                        std__mgr1__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane20_strm1_data        ,
            output  wire                                        mgr1__std__lane20_strm1_data_valid  ,

            // manager 1, lane 21, stream 0      
            input   wire                                        std__mgr1__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane21_strm0_data        ,
            output  wire                                        mgr1__std__lane21_strm0_data_valid  ,

            // manager 1, lane 21, stream 1      
            input   wire                                        std__mgr1__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane21_strm1_data        ,
            output  wire                                        mgr1__std__lane21_strm1_data_valid  ,

            // manager 1, lane 22, stream 0      
            input   wire                                        std__mgr1__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane22_strm0_data        ,
            output  wire                                        mgr1__std__lane22_strm0_data_valid  ,

            // manager 1, lane 22, stream 1      
            input   wire                                        std__mgr1__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane22_strm1_data        ,
            output  wire                                        mgr1__std__lane22_strm1_data_valid  ,

            // manager 1, lane 23, stream 0      
            input   wire                                        std__mgr1__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane23_strm0_data        ,
            output  wire                                        mgr1__std__lane23_strm0_data_valid  ,

            // manager 1, lane 23, stream 1      
            input   wire                                        std__mgr1__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane23_strm1_data        ,
            output  wire                                        mgr1__std__lane23_strm1_data_valid  ,

            // manager 1, lane 24, stream 0      
            input   wire                                        std__mgr1__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane24_strm0_data        ,
            output  wire                                        mgr1__std__lane24_strm0_data_valid  ,

            // manager 1, lane 24, stream 1      
            input   wire                                        std__mgr1__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane24_strm1_data        ,
            output  wire                                        mgr1__std__lane24_strm1_data_valid  ,

            // manager 1, lane 25, stream 0      
            input   wire                                        std__mgr1__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane25_strm0_data        ,
            output  wire                                        mgr1__std__lane25_strm0_data_valid  ,

            // manager 1, lane 25, stream 1      
            input   wire                                        std__mgr1__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane25_strm1_data        ,
            output  wire                                        mgr1__std__lane25_strm1_data_valid  ,

            // manager 1, lane 26, stream 0      
            input   wire                                        std__mgr1__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane26_strm0_data        ,
            output  wire                                        mgr1__std__lane26_strm0_data_valid  ,

            // manager 1, lane 26, stream 1      
            input   wire                                        std__mgr1__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane26_strm1_data        ,
            output  wire                                        mgr1__std__lane26_strm1_data_valid  ,

            // manager 1, lane 27, stream 0      
            input   wire                                        std__mgr1__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane27_strm0_data        ,
            output  wire                                        mgr1__std__lane27_strm0_data_valid  ,

            // manager 1, lane 27, stream 1      
            input   wire                                        std__mgr1__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane27_strm1_data        ,
            output  wire                                        mgr1__std__lane27_strm1_data_valid  ,

            // manager 1, lane 28, stream 0      
            input   wire                                        std__mgr1__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane28_strm0_data        ,
            output  wire                                        mgr1__std__lane28_strm0_data_valid  ,

            // manager 1, lane 28, stream 1      
            input   wire                                        std__mgr1__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane28_strm1_data        ,
            output  wire                                        mgr1__std__lane28_strm1_data_valid  ,

            // manager 1, lane 29, stream 0      
            input   wire                                        std__mgr1__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane29_strm0_data        ,
            output  wire                                        mgr1__std__lane29_strm0_data_valid  ,

            // manager 1, lane 29, stream 1      
            input   wire                                        std__mgr1__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane29_strm1_data        ,
            output  wire                                        mgr1__std__lane29_strm1_data_valid  ,

            // manager 1, lane 30, stream 0      
            input   wire                                        std__mgr1__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane30_strm0_data        ,
            output  wire                                        mgr1__std__lane30_strm0_data_valid  ,

            // manager 1, lane 30, stream 1      
            input   wire                                        std__mgr1__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane30_strm1_data        ,
            output  wire                                        mgr1__std__lane30_strm1_data_valid  ,

            // manager 1, lane 31, stream 0      
            input   wire                                        std__mgr1__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane31_strm0_data        ,
            output  wire                                        mgr1__std__lane31_strm0_data_valid  ,

            // manager 1, lane 31, stream 1      
            input   wire                                        std__mgr1__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr1__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr1__std__lane31_strm1_data        ,
            output  wire                                        mgr1__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 2, lane 0, stream 0      
            input   wire                                        std__mgr2__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane0_strm0_data        ,
            output  wire                                        mgr2__std__lane0_strm0_data_valid  ,

            // manager 2, lane 0, stream 1      
            input   wire                                        std__mgr2__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane0_strm1_data        ,
            output  wire                                        mgr2__std__lane0_strm1_data_valid  ,

            // manager 2, lane 1, stream 0      
            input   wire                                        std__mgr2__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane1_strm0_data        ,
            output  wire                                        mgr2__std__lane1_strm0_data_valid  ,

            // manager 2, lane 1, stream 1      
            input   wire                                        std__mgr2__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane1_strm1_data        ,
            output  wire                                        mgr2__std__lane1_strm1_data_valid  ,

            // manager 2, lane 2, stream 0      
            input   wire                                        std__mgr2__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane2_strm0_data        ,
            output  wire                                        mgr2__std__lane2_strm0_data_valid  ,

            // manager 2, lane 2, stream 1      
            input   wire                                        std__mgr2__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane2_strm1_data        ,
            output  wire                                        mgr2__std__lane2_strm1_data_valid  ,

            // manager 2, lane 3, stream 0      
            input   wire                                        std__mgr2__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane3_strm0_data        ,
            output  wire                                        mgr2__std__lane3_strm0_data_valid  ,

            // manager 2, lane 3, stream 1      
            input   wire                                        std__mgr2__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane3_strm1_data        ,
            output  wire                                        mgr2__std__lane3_strm1_data_valid  ,

            // manager 2, lane 4, stream 0      
            input   wire                                        std__mgr2__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane4_strm0_data        ,
            output  wire                                        mgr2__std__lane4_strm0_data_valid  ,

            // manager 2, lane 4, stream 1      
            input   wire                                        std__mgr2__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane4_strm1_data        ,
            output  wire                                        mgr2__std__lane4_strm1_data_valid  ,

            // manager 2, lane 5, stream 0      
            input   wire                                        std__mgr2__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane5_strm0_data        ,
            output  wire                                        mgr2__std__lane5_strm0_data_valid  ,

            // manager 2, lane 5, stream 1      
            input   wire                                        std__mgr2__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane5_strm1_data        ,
            output  wire                                        mgr2__std__lane5_strm1_data_valid  ,

            // manager 2, lane 6, stream 0      
            input   wire                                        std__mgr2__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane6_strm0_data        ,
            output  wire                                        mgr2__std__lane6_strm0_data_valid  ,

            // manager 2, lane 6, stream 1      
            input   wire                                        std__mgr2__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane6_strm1_data        ,
            output  wire                                        mgr2__std__lane6_strm1_data_valid  ,

            // manager 2, lane 7, stream 0      
            input   wire                                        std__mgr2__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane7_strm0_data        ,
            output  wire                                        mgr2__std__lane7_strm0_data_valid  ,

            // manager 2, lane 7, stream 1      
            input   wire                                        std__mgr2__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane7_strm1_data        ,
            output  wire                                        mgr2__std__lane7_strm1_data_valid  ,

            // manager 2, lane 8, stream 0      
            input   wire                                        std__mgr2__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane8_strm0_data        ,
            output  wire                                        mgr2__std__lane8_strm0_data_valid  ,

            // manager 2, lane 8, stream 1      
            input   wire                                        std__mgr2__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane8_strm1_data        ,
            output  wire                                        mgr2__std__lane8_strm1_data_valid  ,

            // manager 2, lane 9, stream 0      
            input   wire                                        std__mgr2__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane9_strm0_data        ,
            output  wire                                        mgr2__std__lane9_strm0_data_valid  ,

            // manager 2, lane 9, stream 1      
            input   wire                                        std__mgr2__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane9_strm1_data        ,
            output  wire                                        mgr2__std__lane9_strm1_data_valid  ,

            // manager 2, lane 10, stream 0      
            input   wire                                        std__mgr2__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane10_strm0_data        ,
            output  wire                                        mgr2__std__lane10_strm0_data_valid  ,

            // manager 2, lane 10, stream 1      
            input   wire                                        std__mgr2__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane10_strm1_data        ,
            output  wire                                        mgr2__std__lane10_strm1_data_valid  ,

            // manager 2, lane 11, stream 0      
            input   wire                                        std__mgr2__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane11_strm0_data        ,
            output  wire                                        mgr2__std__lane11_strm0_data_valid  ,

            // manager 2, lane 11, stream 1      
            input   wire                                        std__mgr2__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane11_strm1_data        ,
            output  wire                                        mgr2__std__lane11_strm1_data_valid  ,

            // manager 2, lane 12, stream 0      
            input   wire                                        std__mgr2__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane12_strm0_data        ,
            output  wire                                        mgr2__std__lane12_strm0_data_valid  ,

            // manager 2, lane 12, stream 1      
            input   wire                                        std__mgr2__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane12_strm1_data        ,
            output  wire                                        mgr2__std__lane12_strm1_data_valid  ,

            // manager 2, lane 13, stream 0      
            input   wire                                        std__mgr2__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane13_strm0_data        ,
            output  wire                                        mgr2__std__lane13_strm0_data_valid  ,

            // manager 2, lane 13, stream 1      
            input   wire                                        std__mgr2__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane13_strm1_data        ,
            output  wire                                        mgr2__std__lane13_strm1_data_valid  ,

            // manager 2, lane 14, stream 0      
            input   wire                                        std__mgr2__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane14_strm0_data        ,
            output  wire                                        mgr2__std__lane14_strm0_data_valid  ,

            // manager 2, lane 14, stream 1      
            input   wire                                        std__mgr2__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane14_strm1_data        ,
            output  wire                                        mgr2__std__lane14_strm1_data_valid  ,

            // manager 2, lane 15, stream 0      
            input   wire                                        std__mgr2__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane15_strm0_data        ,
            output  wire                                        mgr2__std__lane15_strm0_data_valid  ,

            // manager 2, lane 15, stream 1      
            input   wire                                        std__mgr2__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane15_strm1_data        ,
            output  wire                                        mgr2__std__lane15_strm1_data_valid  ,

            // manager 2, lane 16, stream 0      
            input   wire                                        std__mgr2__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane16_strm0_data        ,
            output  wire                                        mgr2__std__lane16_strm0_data_valid  ,

            // manager 2, lane 16, stream 1      
            input   wire                                        std__mgr2__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane16_strm1_data        ,
            output  wire                                        mgr2__std__lane16_strm1_data_valid  ,

            // manager 2, lane 17, stream 0      
            input   wire                                        std__mgr2__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane17_strm0_data        ,
            output  wire                                        mgr2__std__lane17_strm0_data_valid  ,

            // manager 2, lane 17, stream 1      
            input   wire                                        std__mgr2__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane17_strm1_data        ,
            output  wire                                        mgr2__std__lane17_strm1_data_valid  ,

            // manager 2, lane 18, stream 0      
            input   wire                                        std__mgr2__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane18_strm0_data        ,
            output  wire                                        mgr2__std__lane18_strm0_data_valid  ,

            // manager 2, lane 18, stream 1      
            input   wire                                        std__mgr2__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane18_strm1_data        ,
            output  wire                                        mgr2__std__lane18_strm1_data_valid  ,

            // manager 2, lane 19, stream 0      
            input   wire                                        std__mgr2__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane19_strm0_data        ,
            output  wire                                        mgr2__std__lane19_strm0_data_valid  ,

            // manager 2, lane 19, stream 1      
            input   wire                                        std__mgr2__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane19_strm1_data        ,
            output  wire                                        mgr2__std__lane19_strm1_data_valid  ,

            // manager 2, lane 20, stream 0      
            input   wire                                        std__mgr2__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane20_strm0_data        ,
            output  wire                                        mgr2__std__lane20_strm0_data_valid  ,

            // manager 2, lane 20, stream 1      
            input   wire                                        std__mgr2__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane20_strm1_data        ,
            output  wire                                        mgr2__std__lane20_strm1_data_valid  ,

            // manager 2, lane 21, stream 0      
            input   wire                                        std__mgr2__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane21_strm0_data        ,
            output  wire                                        mgr2__std__lane21_strm0_data_valid  ,

            // manager 2, lane 21, stream 1      
            input   wire                                        std__mgr2__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane21_strm1_data        ,
            output  wire                                        mgr2__std__lane21_strm1_data_valid  ,

            // manager 2, lane 22, stream 0      
            input   wire                                        std__mgr2__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane22_strm0_data        ,
            output  wire                                        mgr2__std__lane22_strm0_data_valid  ,

            // manager 2, lane 22, stream 1      
            input   wire                                        std__mgr2__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane22_strm1_data        ,
            output  wire                                        mgr2__std__lane22_strm1_data_valid  ,

            // manager 2, lane 23, stream 0      
            input   wire                                        std__mgr2__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane23_strm0_data        ,
            output  wire                                        mgr2__std__lane23_strm0_data_valid  ,

            // manager 2, lane 23, stream 1      
            input   wire                                        std__mgr2__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane23_strm1_data        ,
            output  wire                                        mgr2__std__lane23_strm1_data_valid  ,

            // manager 2, lane 24, stream 0      
            input   wire                                        std__mgr2__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane24_strm0_data        ,
            output  wire                                        mgr2__std__lane24_strm0_data_valid  ,

            // manager 2, lane 24, stream 1      
            input   wire                                        std__mgr2__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane24_strm1_data        ,
            output  wire                                        mgr2__std__lane24_strm1_data_valid  ,

            // manager 2, lane 25, stream 0      
            input   wire                                        std__mgr2__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane25_strm0_data        ,
            output  wire                                        mgr2__std__lane25_strm0_data_valid  ,

            // manager 2, lane 25, stream 1      
            input   wire                                        std__mgr2__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane25_strm1_data        ,
            output  wire                                        mgr2__std__lane25_strm1_data_valid  ,

            // manager 2, lane 26, stream 0      
            input   wire                                        std__mgr2__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane26_strm0_data        ,
            output  wire                                        mgr2__std__lane26_strm0_data_valid  ,

            // manager 2, lane 26, stream 1      
            input   wire                                        std__mgr2__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane26_strm1_data        ,
            output  wire                                        mgr2__std__lane26_strm1_data_valid  ,

            // manager 2, lane 27, stream 0      
            input   wire                                        std__mgr2__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane27_strm0_data        ,
            output  wire                                        mgr2__std__lane27_strm0_data_valid  ,

            // manager 2, lane 27, stream 1      
            input   wire                                        std__mgr2__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane27_strm1_data        ,
            output  wire                                        mgr2__std__lane27_strm1_data_valid  ,

            // manager 2, lane 28, stream 0      
            input   wire                                        std__mgr2__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane28_strm0_data        ,
            output  wire                                        mgr2__std__lane28_strm0_data_valid  ,

            // manager 2, lane 28, stream 1      
            input   wire                                        std__mgr2__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane28_strm1_data        ,
            output  wire                                        mgr2__std__lane28_strm1_data_valid  ,

            // manager 2, lane 29, stream 0      
            input   wire                                        std__mgr2__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane29_strm0_data        ,
            output  wire                                        mgr2__std__lane29_strm0_data_valid  ,

            // manager 2, lane 29, stream 1      
            input   wire                                        std__mgr2__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane29_strm1_data        ,
            output  wire                                        mgr2__std__lane29_strm1_data_valid  ,

            // manager 2, lane 30, stream 0      
            input   wire                                        std__mgr2__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane30_strm0_data        ,
            output  wire                                        mgr2__std__lane30_strm0_data_valid  ,

            // manager 2, lane 30, stream 1      
            input   wire                                        std__mgr2__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane30_strm1_data        ,
            output  wire                                        mgr2__std__lane30_strm1_data_valid  ,

            // manager 2, lane 31, stream 0      
            input   wire                                        std__mgr2__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane31_strm0_data        ,
            output  wire                                        mgr2__std__lane31_strm0_data_valid  ,

            // manager 2, lane 31, stream 1      
            input   wire                                        std__mgr2__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr2__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr2__std__lane31_strm1_data        ,
            output  wire                                        mgr2__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 3, lane 0, stream 0      
            input   wire                                        std__mgr3__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane0_strm0_data        ,
            output  wire                                        mgr3__std__lane0_strm0_data_valid  ,

            // manager 3, lane 0, stream 1      
            input   wire                                        std__mgr3__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane0_strm1_data        ,
            output  wire                                        mgr3__std__lane0_strm1_data_valid  ,

            // manager 3, lane 1, stream 0      
            input   wire                                        std__mgr3__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane1_strm0_data        ,
            output  wire                                        mgr3__std__lane1_strm0_data_valid  ,

            // manager 3, lane 1, stream 1      
            input   wire                                        std__mgr3__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane1_strm1_data        ,
            output  wire                                        mgr3__std__lane1_strm1_data_valid  ,

            // manager 3, lane 2, stream 0      
            input   wire                                        std__mgr3__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane2_strm0_data        ,
            output  wire                                        mgr3__std__lane2_strm0_data_valid  ,

            // manager 3, lane 2, stream 1      
            input   wire                                        std__mgr3__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane2_strm1_data        ,
            output  wire                                        mgr3__std__lane2_strm1_data_valid  ,

            // manager 3, lane 3, stream 0      
            input   wire                                        std__mgr3__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane3_strm0_data        ,
            output  wire                                        mgr3__std__lane3_strm0_data_valid  ,

            // manager 3, lane 3, stream 1      
            input   wire                                        std__mgr3__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane3_strm1_data        ,
            output  wire                                        mgr3__std__lane3_strm1_data_valid  ,

            // manager 3, lane 4, stream 0      
            input   wire                                        std__mgr3__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane4_strm0_data        ,
            output  wire                                        mgr3__std__lane4_strm0_data_valid  ,

            // manager 3, lane 4, stream 1      
            input   wire                                        std__mgr3__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane4_strm1_data        ,
            output  wire                                        mgr3__std__lane4_strm1_data_valid  ,

            // manager 3, lane 5, stream 0      
            input   wire                                        std__mgr3__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane5_strm0_data        ,
            output  wire                                        mgr3__std__lane5_strm0_data_valid  ,

            // manager 3, lane 5, stream 1      
            input   wire                                        std__mgr3__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane5_strm1_data        ,
            output  wire                                        mgr3__std__lane5_strm1_data_valid  ,

            // manager 3, lane 6, stream 0      
            input   wire                                        std__mgr3__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane6_strm0_data        ,
            output  wire                                        mgr3__std__lane6_strm0_data_valid  ,

            // manager 3, lane 6, stream 1      
            input   wire                                        std__mgr3__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane6_strm1_data        ,
            output  wire                                        mgr3__std__lane6_strm1_data_valid  ,

            // manager 3, lane 7, stream 0      
            input   wire                                        std__mgr3__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane7_strm0_data        ,
            output  wire                                        mgr3__std__lane7_strm0_data_valid  ,

            // manager 3, lane 7, stream 1      
            input   wire                                        std__mgr3__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane7_strm1_data        ,
            output  wire                                        mgr3__std__lane7_strm1_data_valid  ,

            // manager 3, lane 8, stream 0      
            input   wire                                        std__mgr3__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane8_strm0_data        ,
            output  wire                                        mgr3__std__lane8_strm0_data_valid  ,

            // manager 3, lane 8, stream 1      
            input   wire                                        std__mgr3__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane8_strm1_data        ,
            output  wire                                        mgr3__std__lane8_strm1_data_valid  ,

            // manager 3, lane 9, stream 0      
            input   wire                                        std__mgr3__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane9_strm0_data        ,
            output  wire                                        mgr3__std__lane9_strm0_data_valid  ,

            // manager 3, lane 9, stream 1      
            input   wire                                        std__mgr3__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane9_strm1_data        ,
            output  wire                                        mgr3__std__lane9_strm1_data_valid  ,

            // manager 3, lane 10, stream 0      
            input   wire                                        std__mgr3__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane10_strm0_data        ,
            output  wire                                        mgr3__std__lane10_strm0_data_valid  ,

            // manager 3, lane 10, stream 1      
            input   wire                                        std__mgr3__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane10_strm1_data        ,
            output  wire                                        mgr3__std__lane10_strm1_data_valid  ,

            // manager 3, lane 11, stream 0      
            input   wire                                        std__mgr3__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane11_strm0_data        ,
            output  wire                                        mgr3__std__lane11_strm0_data_valid  ,

            // manager 3, lane 11, stream 1      
            input   wire                                        std__mgr3__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane11_strm1_data        ,
            output  wire                                        mgr3__std__lane11_strm1_data_valid  ,

            // manager 3, lane 12, stream 0      
            input   wire                                        std__mgr3__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane12_strm0_data        ,
            output  wire                                        mgr3__std__lane12_strm0_data_valid  ,

            // manager 3, lane 12, stream 1      
            input   wire                                        std__mgr3__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane12_strm1_data        ,
            output  wire                                        mgr3__std__lane12_strm1_data_valid  ,

            // manager 3, lane 13, stream 0      
            input   wire                                        std__mgr3__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane13_strm0_data        ,
            output  wire                                        mgr3__std__lane13_strm0_data_valid  ,

            // manager 3, lane 13, stream 1      
            input   wire                                        std__mgr3__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane13_strm1_data        ,
            output  wire                                        mgr3__std__lane13_strm1_data_valid  ,

            // manager 3, lane 14, stream 0      
            input   wire                                        std__mgr3__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane14_strm0_data        ,
            output  wire                                        mgr3__std__lane14_strm0_data_valid  ,

            // manager 3, lane 14, stream 1      
            input   wire                                        std__mgr3__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane14_strm1_data        ,
            output  wire                                        mgr3__std__lane14_strm1_data_valid  ,

            // manager 3, lane 15, stream 0      
            input   wire                                        std__mgr3__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane15_strm0_data        ,
            output  wire                                        mgr3__std__lane15_strm0_data_valid  ,

            // manager 3, lane 15, stream 1      
            input   wire                                        std__mgr3__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane15_strm1_data        ,
            output  wire                                        mgr3__std__lane15_strm1_data_valid  ,

            // manager 3, lane 16, stream 0      
            input   wire                                        std__mgr3__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane16_strm0_data        ,
            output  wire                                        mgr3__std__lane16_strm0_data_valid  ,

            // manager 3, lane 16, stream 1      
            input   wire                                        std__mgr3__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane16_strm1_data        ,
            output  wire                                        mgr3__std__lane16_strm1_data_valid  ,

            // manager 3, lane 17, stream 0      
            input   wire                                        std__mgr3__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane17_strm0_data        ,
            output  wire                                        mgr3__std__lane17_strm0_data_valid  ,

            // manager 3, lane 17, stream 1      
            input   wire                                        std__mgr3__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane17_strm1_data        ,
            output  wire                                        mgr3__std__lane17_strm1_data_valid  ,

            // manager 3, lane 18, stream 0      
            input   wire                                        std__mgr3__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane18_strm0_data        ,
            output  wire                                        mgr3__std__lane18_strm0_data_valid  ,

            // manager 3, lane 18, stream 1      
            input   wire                                        std__mgr3__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane18_strm1_data        ,
            output  wire                                        mgr3__std__lane18_strm1_data_valid  ,

            // manager 3, lane 19, stream 0      
            input   wire                                        std__mgr3__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane19_strm0_data        ,
            output  wire                                        mgr3__std__lane19_strm0_data_valid  ,

            // manager 3, lane 19, stream 1      
            input   wire                                        std__mgr3__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane19_strm1_data        ,
            output  wire                                        mgr3__std__lane19_strm1_data_valid  ,

            // manager 3, lane 20, stream 0      
            input   wire                                        std__mgr3__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane20_strm0_data        ,
            output  wire                                        mgr3__std__lane20_strm0_data_valid  ,

            // manager 3, lane 20, stream 1      
            input   wire                                        std__mgr3__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane20_strm1_data        ,
            output  wire                                        mgr3__std__lane20_strm1_data_valid  ,

            // manager 3, lane 21, stream 0      
            input   wire                                        std__mgr3__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane21_strm0_data        ,
            output  wire                                        mgr3__std__lane21_strm0_data_valid  ,

            // manager 3, lane 21, stream 1      
            input   wire                                        std__mgr3__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane21_strm1_data        ,
            output  wire                                        mgr3__std__lane21_strm1_data_valid  ,

            // manager 3, lane 22, stream 0      
            input   wire                                        std__mgr3__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane22_strm0_data        ,
            output  wire                                        mgr3__std__lane22_strm0_data_valid  ,

            // manager 3, lane 22, stream 1      
            input   wire                                        std__mgr3__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane22_strm1_data        ,
            output  wire                                        mgr3__std__lane22_strm1_data_valid  ,

            // manager 3, lane 23, stream 0      
            input   wire                                        std__mgr3__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane23_strm0_data        ,
            output  wire                                        mgr3__std__lane23_strm0_data_valid  ,

            // manager 3, lane 23, stream 1      
            input   wire                                        std__mgr3__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane23_strm1_data        ,
            output  wire                                        mgr3__std__lane23_strm1_data_valid  ,

            // manager 3, lane 24, stream 0      
            input   wire                                        std__mgr3__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane24_strm0_data        ,
            output  wire                                        mgr3__std__lane24_strm0_data_valid  ,

            // manager 3, lane 24, stream 1      
            input   wire                                        std__mgr3__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane24_strm1_data        ,
            output  wire                                        mgr3__std__lane24_strm1_data_valid  ,

            // manager 3, lane 25, stream 0      
            input   wire                                        std__mgr3__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane25_strm0_data        ,
            output  wire                                        mgr3__std__lane25_strm0_data_valid  ,

            // manager 3, lane 25, stream 1      
            input   wire                                        std__mgr3__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane25_strm1_data        ,
            output  wire                                        mgr3__std__lane25_strm1_data_valid  ,

            // manager 3, lane 26, stream 0      
            input   wire                                        std__mgr3__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane26_strm0_data        ,
            output  wire                                        mgr3__std__lane26_strm0_data_valid  ,

            // manager 3, lane 26, stream 1      
            input   wire                                        std__mgr3__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane26_strm1_data        ,
            output  wire                                        mgr3__std__lane26_strm1_data_valid  ,

            // manager 3, lane 27, stream 0      
            input   wire                                        std__mgr3__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane27_strm0_data        ,
            output  wire                                        mgr3__std__lane27_strm0_data_valid  ,

            // manager 3, lane 27, stream 1      
            input   wire                                        std__mgr3__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane27_strm1_data        ,
            output  wire                                        mgr3__std__lane27_strm1_data_valid  ,

            // manager 3, lane 28, stream 0      
            input   wire                                        std__mgr3__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane28_strm0_data        ,
            output  wire                                        mgr3__std__lane28_strm0_data_valid  ,

            // manager 3, lane 28, stream 1      
            input   wire                                        std__mgr3__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane28_strm1_data        ,
            output  wire                                        mgr3__std__lane28_strm1_data_valid  ,

            // manager 3, lane 29, stream 0      
            input   wire                                        std__mgr3__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane29_strm0_data        ,
            output  wire                                        mgr3__std__lane29_strm0_data_valid  ,

            // manager 3, lane 29, stream 1      
            input   wire                                        std__mgr3__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane29_strm1_data        ,
            output  wire                                        mgr3__std__lane29_strm1_data_valid  ,

            // manager 3, lane 30, stream 0      
            input   wire                                        std__mgr3__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane30_strm0_data        ,
            output  wire                                        mgr3__std__lane30_strm0_data_valid  ,

            // manager 3, lane 30, stream 1      
            input   wire                                        std__mgr3__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane30_strm1_data        ,
            output  wire                                        mgr3__std__lane30_strm1_data_valid  ,

            // manager 3, lane 31, stream 0      
            input   wire                                        std__mgr3__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane31_strm0_data        ,
            output  wire                                        mgr3__std__lane31_strm0_data_valid  ,

            // manager 3, lane 31, stream 1      
            input   wire                                        std__mgr3__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr3__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr3__std__lane31_strm1_data        ,
            output  wire                                        mgr3__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 4, lane 0, stream 0      
            input   wire                                        std__mgr4__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane0_strm0_data        ,
            output  wire                                        mgr4__std__lane0_strm0_data_valid  ,

            // manager 4, lane 0, stream 1      
            input   wire                                        std__mgr4__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane0_strm1_data        ,
            output  wire                                        mgr4__std__lane0_strm1_data_valid  ,

            // manager 4, lane 1, stream 0      
            input   wire                                        std__mgr4__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane1_strm0_data        ,
            output  wire                                        mgr4__std__lane1_strm0_data_valid  ,

            // manager 4, lane 1, stream 1      
            input   wire                                        std__mgr4__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane1_strm1_data        ,
            output  wire                                        mgr4__std__lane1_strm1_data_valid  ,

            // manager 4, lane 2, stream 0      
            input   wire                                        std__mgr4__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane2_strm0_data        ,
            output  wire                                        mgr4__std__lane2_strm0_data_valid  ,

            // manager 4, lane 2, stream 1      
            input   wire                                        std__mgr4__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane2_strm1_data        ,
            output  wire                                        mgr4__std__lane2_strm1_data_valid  ,

            // manager 4, lane 3, stream 0      
            input   wire                                        std__mgr4__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane3_strm0_data        ,
            output  wire                                        mgr4__std__lane3_strm0_data_valid  ,

            // manager 4, lane 3, stream 1      
            input   wire                                        std__mgr4__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane3_strm1_data        ,
            output  wire                                        mgr4__std__lane3_strm1_data_valid  ,

            // manager 4, lane 4, stream 0      
            input   wire                                        std__mgr4__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane4_strm0_data        ,
            output  wire                                        mgr4__std__lane4_strm0_data_valid  ,

            // manager 4, lane 4, stream 1      
            input   wire                                        std__mgr4__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane4_strm1_data        ,
            output  wire                                        mgr4__std__lane4_strm1_data_valid  ,

            // manager 4, lane 5, stream 0      
            input   wire                                        std__mgr4__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane5_strm0_data        ,
            output  wire                                        mgr4__std__lane5_strm0_data_valid  ,

            // manager 4, lane 5, stream 1      
            input   wire                                        std__mgr4__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane5_strm1_data        ,
            output  wire                                        mgr4__std__lane5_strm1_data_valid  ,

            // manager 4, lane 6, stream 0      
            input   wire                                        std__mgr4__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane6_strm0_data        ,
            output  wire                                        mgr4__std__lane6_strm0_data_valid  ,

            // manager 4, lane 6, stream 1      
            input   wire                                        std__mgr4__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane6_strm1_data        ,
            output  wire                                        mgr4__std__lane6_strm1_data_valid  ,

            // manager 4, lane 7, stream 0      
            input   wire                                        std__mgr4__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane7_strm0_data        ,
            output  wire                                        mgr4__std__lane7_strm0_data_valid  ,

            // manager 4, lane 7, stream 1      
            input   wire                                        std__mgr4__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane7_strm1_data        ,
            output  wire                                        mgr4__std__lane7_strm1_data_valid  ,

            // manager 4, lane 8, stream 0      
            input   wire                                        std__mgr4__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane8_strm0_data        ,
            output  wire                                        mgr4__std__lane8_strm0_data_valid  ,

            // manager 4, lane 8, stream 1      
            input   wire                                        std__mgr4__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane8_strm1_data        ,
            output  wire                                        mgr4__std__lane8_strm1_data_valid  ,

            // manager 4, lane 9, stream 0      
            input   wire                                        std__mgr4__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane9_strm0_data        ,
            output  wire                                        mgr4__std__lane9_strm0_data_valid  ,

            // manager 4, lane 9, stream 1      
            input   wire                                        std__mgr4__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane9_strm1_data        ,
            output  wire                                        mgr4__std__lane9_strm1_data_valid  ,

            // manager 4, lane 10, stream 0      
            input   wire                                        std__mgr4__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane10_strm0_data        ,
            output  wire                                        mgr4__std__lane10_strm0_data_valid  ,

            // manager 4, lane 10, stream 1      
            input   wire                                        std__mgr4__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane10_strm1_data        ,
            output  wire                                        mgr4__std__lane10_strm1_data_valid  ,

            // manager 4, lane 11, stream 0      
            input   wire                                        std__mgr4__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane11_strm0_data        ,
            output  wire                                        mgr4__std__lane11_strm0_data_valid  ,

            // manager 4, lane 11, stream 1      
            input   wire                                        std__mgr4__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane11_strm1_data        ,
            output  wire                                        mgr4__std__lane11_strm1_data_valid  ,

            // manager 4, lane 12, stream 0      
            input   wire                                        std__mgr4__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane12_strm0_data        ,
            output  wire                                        mgr4__std__lane12_strm0_data_valid  ,

            // manager 4, lane 12, stream 1      
            input   wire                                        std__mgr4__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane12_strm1_data        ,
            output  wire                                        mgr4__std__lane12_strm1_data_valid  ,

            // manager 4, lane 13, stream 0      
            input   wire                                        std__mgr4__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane13_strm0_data        ,
            output  wire                                        mgr4__std__lane13_strm0_data_valid  ,

            // manager 4, lane 13, stream 1      
            input   wire                                        std__mgr4__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane13_strm1_data        ,
            output  wire                                        mgr4__std__lane13_strm1_data_valid  ,

            // manager 4, lane 14, stream 0      
            input   wire                                        std__mgr4__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane14_strm0_data        ,
            output  wire                                        mgr4__std__lane14_strm0_data_valid  ,

            // manager 4, lane 14, stream 1      
            input   wire                                        std__mgr4__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane14_strm1_data        ,
            output  wire                                        mgr4__std__lane14_strm1_data_valid  ,

            // manager 4, lane 15, stream 0      
            input   wire                                        std__mgr4__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane15_strm0_data        ,
            output  wire                                        mgr4__std__lane15_strm0_data_valid  ,

            // manager 4, lane 15, stream 1      
            input   wire                                        std__mgr4__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane15_strm1_data        ,
            output  wire                                        mgr4__std__lane15_strm1_data_valid  ,

            // manager 4, lane 16, stream 0      
            input   wire                                        std__mgr4__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane16_strm0_data        ,
            output  wire                                        mgr4__std__lane16_strm0_data_valid  ,

            // manager 4, lane 16, stream 1      
            input   wire                                        std__mgr4__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane16_strm1_data        ,
            output  wire                                        mgr4__std__lane16_strm1_data_valid  ,

            // manager 4, lane 17, stream 0      
            input   wire                                        std__mgr4__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane17_strm0_data        ,
            output  wire                                        mgr4__std__lane17_strm0_data_valid  ,

            // manager 4, lane 17, stream 1      
            input   wire                                        std__mgr4__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane17_strm1_data        ,
            output  wire                                        mgr4__std__lane17_strm1_data_valid  ,

            // manager 4, lane 18, stream 0      
            input   wire                                        std__mgr4__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane18_strm0_data        ,
            output  wire                                        mgr4__std__lane18_strm0_data_valid  ,

            // manager 4, lane 18, stream 1      
            input   wire                                        std__mgr4__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane18_strm1_data        ,
            output  wire                                        mgr4__std__lane18_strm1_data_valid  ,

            // manager 4, lane 19, stream 0      
            input   wire                                        std__mgr4__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane19_strm0_data        ,
            output  wire                                        mgr4__std__lane19_strm0_data_valid  ,

            // manager 4, lane 19, stream 1      
            input   wire                                        std__mgr4__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane19_strm1_data        ,
            output  wire                                        mgr4__std__lane19_strm1_data_valid  ,

            // manager 4, lane 20, stream 0      
            input   wire                                        std__mgr4__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane20_strm0_data        ,
            output  wire                                        mgr4__std__lane20_strm0_data_valid  ,

            // manager 4, lane 20, stream 1      
            input   wire                                        std__mgr4__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane20_strm1_data        ,
            output  wire                                        mgr4__std__lane20_strm1_data_valid  ,

            // manager 4, lane 21, stream 0      
            input   wire                                        std__mgr4__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane21_strm0_data        ,
            output  wire                                        mgr4__std__lane21_strm0_data_valid  ,

            // manager 4, lane 21, stream 1      
            input   wire                                        std__mgr4__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane21_strm1_data        ,
            output  wire                                        mgr4__std__lane21_strm1_data_valid  ,

            // manager 4, lane 22, stream 0      
            input   wire                                        std__mgr4__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane22_strm0_data        ,
            output  wire                                        mgr4__std__lane22_strm0_data_valid  ,

            // manager 4, lane 22, stream 1      
            input   wire                                        std__mgr4__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane22_strm1_data        ,
            output  wire                                        mgr4__std__lane22_strm1_data_valid  ,

            // manager 4, lane 23, stream 0      
            input   wire                                        std__mgr4__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane23_strm0_data        ,
            output  wire                                        mgr4__std__lane23_strm0_data_valid  ,

            // manager 4, lane 23, stream 1      
            input   wire                                        std__mgr4__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane23_strm1_data        ,
            output  wire                                        mgr4__std__lane23_strm1_data_valid  ,

            // manager 4, lane 24, stream 0      
            input   wire                                        std__mgr4__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane24_strm0_data        ,
            output  wire                                        mgr4__std__lane24_strm0_data_valid  ,

            // manager 4, lane 24, stream 1      
            input   wire                                        std__mgr4__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane24_strm1_data        ,
            output  wire                                        mgr4__std__lane24_strm1_data_valid  ,

            // manager 4, lane 25, stream 0      
            input   wire                                        std__mgr4__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane25_strm0_data        ,
            output  wire                                        mgr4__std__lane25_strm0_data_valid  ,

            // manager 4, lane 25, stream 1      
            input   wire                                        std__mgr4__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane25_strm1_data        ,
            output  wire                                        mgr4__std__lane25_strm1_data_valid  ,

            // manager 4, lane 26, stream 0      
            input   wire                                        std__mgr4__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane26_strm0_data        ,
            output  wire                                        mgr4__std__lane26_strm0_data_valid  ,

            // manager 4, lane 26, stream 1      
            input   wire                                        std__mgr4__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane26_strm1_data        ,
            output  wire                                        mgr4__std__lane26_strm1_data_valid  ,

            // manager 4, lane 27, stream 0      
            input   wire                                        std__mgr4__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane27_strm0_data        ,
            output  wire                                        mgr4__std__lane27_strm0_data_valid  ,

            // manager 4, lane 27, stream 1      
            input   wire                                        std__mgr4__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane27_strm1_data        ,
            output  wire                                        mgr4__std__lane27_strm1_data_valid  ,

            // manager 4, lane 28, stream 0      
            input   wire                                        std__mgr4__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane28_strm0_data        ,
            output  wire                                        mgr4__std__lane28_strm0_data_valid  ,

            // manager 4, lane 28, stream 1      
            input   wire                                        std__mgr4__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane28_strm1_data        ,
            output  wire                                        mgr4__std__lane28_strm1_data_valid  ,

            // manager 4, lane 29, stream 0      
            input   wire                                        std__mgr4__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane29_strm0_data        ,
            output  wire                                        mgr4__std__lane29_strm0_data_valid  ,

            // manager 4, lane 29, stream 1      
            input   wire                                        std__mgr4__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane29_strm1_data        ,
            output  wire                                        mgr4__std__lane29_strm1_data_valid  ,

            // manager 4, lane 30, stream 0      
            input   wire                                        std__mgr4__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane30_strm0_data        ,
            output  wire                                        mgr4__std__lane30_strm0_data_valid  ,

            // manager 4, lane 30, stream 1      
            input   wire                                        std__mgr4__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane30_strm1_data        ,
            output  wire                                        mgr4__std__lane30_strm1_data_valid  ,

            // manager 4, lane 31, stream 0      
            input   wire                                        std__mgr4__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane31_strm0_data        ,
            output  wire                                        mgr4__std__lane31_strm0_data_valid  ,

            // manager 4, lane 31, stream 1      
            input   wire                                        std__mgr4__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr4__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr4__std__lane31_strm1_data        ,
            output  wire                                        mgr4__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 5, lane 0, stream 0      
            input   wire                                        std__mgr5__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane0_strm0_data        ,
            output  wire                                        mgr5__std__lane0_strm0_data_valid  ,

            // manager 5, lane 0, stream 1      
            input   wire                                        std__mgr5__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane0_strm1_data        ,
            output  wire                                        mgr5__std__lane0_strm1_data_valid  ,

            // manager 5, lane 1, stream 0      
            input   wire                                        std__mgr5__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane1_strm0_data        ,
            output  wire                                        mgr5__std__lane1_strm0_data_valid  ,

            // manager 5, lane 1, stream 1      
            input   wire                                        std__mgr5__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane1_strm1_data        ,
            output  wire                                        mgr5__std__lane1_strm1_data_valid  ,

            // manager 5, lane 2, stream 0      
            input   wire                                        std__mgr5__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane2_strm0_data        ,
            output  wire                                        mgr5__std__lane2_strm0_data_valid  ,

            // manager 5, lane 2, stream 1      
            input   wire                                        std__mgr5__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane2_strm1_data        ,
            output  wire                                        mgr5__std__lane2_strm1_data_valid  ,

            // manager 5, lane 3, stream 0      
            input   wire                                        std__mgr5__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane3_strm0_data        ,
            output  wire                                        mgr5__std__lane3_strm0_data_valid  ,

            // manager 5, lane 3, stream 1      
            input   wire                                        std__mgr5__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane3_strm1_data        ,
            output  wire                                        mgr5__std__lane3_strm1_data_valid  ,

            // manager 5, lane 4, stream 0      
            input   wire                                        std__mgr5__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane4_strm0_data        ,
            output  wire                                        mgr5__std__lane4_strm0_data_valid  ,

            // manager 5, lane 4, stream 1      
            input   wire                                        std__mgr5__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane4_strm1_data        ,
            output  wire                                        mgr5__std__lane4_strm1_data_valid  ,

            // manager 5, lane 5, stream 0      
            input   wire                                        std__mgr5__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane5_strm0_data        ,
            output  wire                                        mgr5__std__lane5_strm0_data_valid  ,

            // manager 5, lane 5, stream 1      
            input   wire                                        std__mgr5__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane5_strm1_data        ,
            output  wire                                        mgr5__std__lane5_strm1_data_valid  ,

            // manager 5, lane 6, stream 0      
            input   wire                                        std__mgr5__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane6_strm0_data        ,
            output  wire                                        mgr5__std__lane6_strm0_data_valid  ,

            // manager 5, lane 6, stream 1      
            input   wire                                        std__mgr5__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane6_strm1_data        ,
            output  wire                                        mgr5__std__lane6_strm1_data_valid  ,

            // manager 5, lane 7, stream 0      
            input   wire                                        std__mgr5__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane7_strm0_data        ,
            output  wire                                        mgr5__std__lane7_strm0_data_valid  ,

            // manager 5, lane 7, stream 1      
            input   wire                                        std__mgr5__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane7_strm1_data        ,
            output  wire                                        mgr5__std__lane7_strm1_data_valid  ,

            // manager 5, lane 8, stream 0      
            input   wire                                        std__mgr5__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane8_strm0_data        ,
            output  wire                                        mgr5__std__lane8_strm0_data_valid  ,

            // manager 5, lane 8, stream 1      
            input   wire                                        std__mgr5__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane8_strm1_data        ,
            output  wire                                        mgr5__std__lane8_strm1_data_valid  ,

            // manager 5, lane 9, stream 0      
            input   wire                                        std__mgr5__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane9_strm0_data        ,
            output  wire                                        mgr5__std__lane9_strm0_data_valid  ,

            // manager 5, lane 9, stream 1      
            input   wire                                        std__mgr5__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane9_strm1_data        ,
            output  wire                                        mgr5__std__lane9_strm1_data_valid  ,

            // manager 5, lane 10, stream 0      
            input   wire                                        std__mgr5__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane10_strm0_data        ,
            output  wire                                        mgr5__std__lane10_strm0_data_valid  ,

            // manager 5, lane 10, stream 1      
            input   wire                                        std__mgr5__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane10_strm1_data        ,
            output  wire                                        mgr5__std__lane10_strm1_data_valid  ,

            // manager 5, lane 11, stream 0      
            input   wire                                        std__mgr5__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane11_strm0_data        ,
            output  wire                                        mgr5__std__lane11_strm0_data_valid  ,

            // manager 5, lane 11, stream 1      
            input   wire                                        std__mgr5__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane11_strm1_data        ,
            output  wire                                        mgr5__std__lane11_strm1_data_valid  ,

            // manager 5, lane 12, stream 0      
            input   wire                                        std__mgr5__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane12_strm0_data        ,
            output  wire                                        mgr5__std__lane12_strm0_data_valid  ,

            // manager 5, lane 12, stream 1      
            input   wire                                        std__mgr5__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane12_strm1_data        ,
            output  wire                                        mgr5__std__lane12_strm1_data_valid  ,

            // manager 5, lane 13, stream 0      
            input   wire                                        std__mgr5__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane13_strm0_data        ,
            output  wire                                        mgr5__std__lane13_strm0_data_valid  ,

            // manager 5, lane 13, stream 1      
            input   wire                                        std__mgr5__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane13_strm1_data        ,
            output  wire                                        mgr5__std__lane13_strm1_data_valid  ,

            // manager 5, lane 14, stream 0      
            input   wire                                        std__mgr5__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane14_strm0_data        ,
            output  wire                                        mgr5__std__lane14_strm0_data_valid  ,

            // manager 5, lane 14, stream 1      
            input   wire                                        std__mgr5__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane14_strm1_data        ,
            output  wire                                        mgr5__std__lane14_strm1_data_valid  ,

            // manager 5, lane 15, stream 0      
            input   wire                                        std__mgr5__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane15_strm0_data        ,
            output  wire                                        mgr5__std__lane15_strm0_data_valid  ,

            // manager 5, lane 15, stream 1      
            input   wire                                        std__mgr5__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane15_strm1_data        ,
            output  wire                                        mgr5__std__lane15_strm1_data_valid  ,

            // manager 5, lane 16, stream 0      
            input   wire                                        std__mgr5__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane16_strm0_data        ,
            output  wire                                        mgr5__std__lane16_strm0_data_valid  ,

            // manager 5, lane 16, stream 1      
            input   wire                                        std__mgr5__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane16_strm1_data        ,
            output  wire                                        mgr5__std__lane16_strm1_data_valid  ,

            // manager 5, lane 17, stream 0      
            input   wire                                        std__mgr5__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane17_strm0_data        ,
            output  wire                                        mgr5__std__lane17_strm0_data_valid  ,

            // manager 5, lane 17, stream 1      
            input   wire                                        std__mgr5__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane17_strm1_data        ,
            output  wire                                        mgr5__std__lane17_strm1_data_valid  ,

            // manager 5, lane 18, stream 0      
            input   wire                                        std__mgr5__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane18_strm0_data        ,
            output  wire                                        mgr5__std__lane18_strm0_data_valid  ,

            // manager 5, lane 18, stream 1      
            input   wire                                        std__mgr5__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane18_strm1_data        ,
            output  wire                                        mgr5__std__lane18_strm1_data_valid  ,

            // manager 5, lane 19, stream 0      
            input   wire                                        std__mgr5__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane19_strm0_data        ,
            output  wire                                        mgr5__std__lane19_strm0_data_valid  ,

            // manager 5, lane 19, stream 1      
            input   wire                                        std__mgr5__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane19_strm1_data        ,
            output  wire                                        mgr5__std__lane19_strm1_data_valid  ,

            // manager 5, lane 20, stream 0      
            input   wire                                        std__mgr5__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane20_strm0_data        ,
            output  wire                                        mgr5__std__lane20_strm0_data_valid  ,

            // manager 5, lane 20, stream 1      
            input   wire                                        std__mgr5__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane20_strm1_data        ,
            output  wire                                        mgr5__std__lane20_strm1_data_valid  ,

            // manager 5, lane 21, stream 0      
            input   wire                                        std__mgr5__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane21_strm0_data        ,
            output  wire                                        mgr5__std__lane21_strm0_data_valid  ,

            // manager 5, lane 21, stream 1      
            input   wire                                        std__mgr5__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane21_strm1_data        ,
            output  wire                                        mgr5__std__lane21_strm1_data_valid  ,

            // manager 5, lane 22, stream 0      
            input   wire                                        std__mgr5__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane22_strm0_data        ,
            output  wire                                        mgr5__std__lane22_strm0_data_valid  ,

            // manager 5, lane 22, stream 1      
            input   wire                                        std__mgr5__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane22_strm1_data        ,
            output  wire                                        mgr5__std__lane22_strm1_data_valid  ,

            // manager 5, lane 23, stream 0      
            input   wire                                        std__mgr5__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane23_strm0_data        ,
            output  wire                                        mgr5__std__lane23_strm0_data_valid  ,

            // manager 5, lane 23, stream 1      
            input   wire                                        std__mgr5__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane23_strm1_data        ,
            output  wire                                        mgr5__std__lane23_strm1_data_valid  ,

            // manager 5, lane 24, stream 0      
            input   wire                                        std__mgr5__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane24_strm0_data        ,
            output  wire                                        mgr5__std__lane24_strm0_data_valid  ,

            // manager 5, lane 24, stream 1      
            input   wire                                        std__mgr5__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane24_strm1_data        ,
            output  wire                                        mgr5__std__lane24_strm1_data_valid  ,

            // manager 5, lane 25, stream 0      
            input   wire                                        std__mgr5__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane25_strm0_data        ,
            output  wire                                        mgr5__std__lane25_strm0_data_valid  ,

            // manager 5, lane 25, stream 1      
            input   wire                                        std__mgr5__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane25_strm1_data        ,
            output  wire                                        mgr5__std__lane25_strm1_data_valid  ,

            // manager 5, lane 26, stream 0      
            input   wire                                        std__mgr5__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane26_strm0_data        ,
            output  wire                                        mgr5__std__lane26_strm0_data_valid  ,

            // manager 5, lane 26, stream 1      
            input   wire                                        std__mgr5__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane26_strm1_data        ,
            output  wire                                        mgr5__std__lane26_strm1_data_valid  ,

            // manager 5, lane 27, stream 0      
            input   wire                                        std__mgr5__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane27_strm0_data        ,
            output  wire                                        mgr5__std__lane27_strm0_data_valid  ,

            // manager 5, lane 27, stream 1      
            input   wire                                        std__mgr5__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane27_strm1_data        ,
            output  wire                                        mgr5__std__lane27_strm1_data_valid  ,

            // manager 5, lane 28, stream 0      
            input   wire                                        std__mgr5__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane28_strm0_data        ,
            output  wire                                        mgr5__std__lane28_strm0_data_valid  ,

            // manager 5, lane 28, stream 1      
            input   wire                                        std__mgr5__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane28_strm1_data        ,
            output  wire                                        mgr5__std__lane28_strm1_data_valid  ,

            // manager 5, lane 29, stream 0      
            input   wire                                        std__mgr5__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane29_strm0_data        ,
            output  wire                                        mgr5__std__lane29_strm0_data_valid  ,

            // manager 5, lane 29, stream 1      
            input   wire                                        std__mgr5__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane29_strm1_data        ,
            output  wire                                        mgr5__std__lane29_strm1_data_valid  ,

            // manager 5, lane 30, stream 0      
            input   wire                                        std__mgr5__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane30_strm0_data        ,
            output  wire                                        mgr5__std__lane30_strm0_data_valid  ,

            // manager 5, lane 30, stream 1      
            input   wire                                        std__mgr5__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane30_strm1_data        ,
            output  wire                                        mgr5__std__lane30_strm1_data_valid  ,

            // manager 5, lane 31, stream 0      
            input   wire                                        std__mgr5__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane31_strm0_data        ,
            output  wire                                        mgr5__std__lane31_strm0_data_valid  ,

            // manager 5, lane 31, stream 1      
            input   wire                                        std__mgr5__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr5__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr5__std__lane31_strm1_data        ,
            output  wire                                        mgr5__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 6, lane 0, stream 0      
            input   wire                                        std__mgr6__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane0_strm0_data        ,
            output  wire                                        mgr6__std__lane0_strm0_data_valid  ,

            // manager 6, lane 0, stream 1      
            input   wire                                        std__mgr6__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane0_strm1_data        ,
            output  wire                                        mgr6__std__lane0_strm1_data_valid  ,

            // manager 6, lane 1, stream 0      
            input   wire                                        std__mgr6__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane1_strm0_data        ,
            output  wire                                        mgr6__std__lane1_strm0_data_valid  ,

            // manager 6, lane 1, stream 1      
            input   wire                                        std__mgr6__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane1_strm1_data        ,
            output  wire                                        mgr6__std__lane1_strm1_data_valid  ,

            // manager 6, lane 2, stream 0      
            input   wire                                        std__mgr6__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane2_strm0_data        ,
            output  wire                                        mgr6__std__lane2_strm0_data_valid  ,

            // manager 6, lane 2, stream 1      
            input   wire                                        std__mgr6__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane2_strm1_data        ,
            output  wire                                        mgr6__std__lane2_strm1_data_valid  ,

            // manager 6, lane 3, stream 0      
            input   wire                                        std__mgr6__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane3_strm0_data        ,
            output  wire                                        mgr6__std__lane3_strm0_data_valid  ,

            // manager 6, lane 3, stream 1      
            input   wire                                        std__mgr6__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane3_strm1_data        ,
            output  wire                                        mgr6__std__lane3_strm1_data_valid  ,

            // manager 6, lane 4, stream 0      
            input   wire                                        std__mgr6__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane4_strm0_data        ,
            output  wire                                        mgr6__std__lane4_strm0_data_valid  ,

            // manager 6, lane 4, stream 1      
            input   wire                                        std__mgr6__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane4_strm1_data        ,
            output  wire                                        mgr6__std__lane4_strm1_data_valid  ,

            // manager 6, lane 5, stream 0      
            input   wire                                        std__mgr6__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane5_strm0_data        ,
            output  wire                                        mgr6__std__lane5_strm0_data_valid  ,

            // manager 6, lane 5, stream 1      
            input   wire                                        std__mgr6__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane5_strm1_data        ,
            output  wire                                        mgr6__std__lane5_strm1_data_valid  ,

            // manager 6, lane 6, stream 0      
            input   wire                                        std__mgr6__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane6_strm0_data        ,
            output  wire                                        mgr6__std__lane6_strm0_data_valid  ,

            // manager 6, lane 6, stream 1      
            input   wire                                        std__mgr6__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane6_strm1_data        ,
            output  wire                                        mgr6__std__lane6_strm1_data_valid  ,

            // manager 6, lane 7, stream 0      
            input   wire                                        std__mgr6__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane7_strm0_data        ,
            output  wire                                        mgr6__std__lane7_strm0_data_valid  ,

            // manager 6, lane 7, stream 1      
            input   wire                                        std__mgr6__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane7_strm1_data        ,
            output  wire                                        mgr6__std__lane7_strm1_data_valid  ,

            // manager 6, lane 8, stream 0      
            input   wire                                        std__mgr6__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane8_strm0_data        ,
            output  wire                                        mgr6__std__lane8_strm0_data_valid  ,

            // manager 6, lane 8, stream 1      
            input   wire                                        std__mgr6__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane8_strm1_data        ,
            output  wire                                        mgr6__std__lane8_strm1_data_valid  ,

            // manager 6, lane 9, stream 0      
            input   wire                                        std__mgr6__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane9_strm0_data        ,
            output  wire                                        mgr6__std__lane9_strm0_data_valid  ,

            // manager 6, lane 9, stream 1      
            input   wire                                        std__mgr6__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane9_strm1_data        ,
            output  wire                                        mgr6__std__lane9_strm1_data_valid  ,

            // manager 6, lane 10, stream 0      
            input   wire                                        std__mgr6__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane10_strm0_data        ,
            output  wire                                        mgr6__std__lane10_strm0_data_valid  ,

            // manager 6, lane 10, stream 1      
            input   wire                                        std__mgr6__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane10_strm1_data        ,
            output  wire                                        mgr6__std__lane10_strm1_data_valid  ,

            // manager 6, lane 11, stream 0      
            input   wire                                        std__mgr6__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane11_strm0_data        ,
            output  wire                                        mgr6__std__lane11_strm0_data_valid  ,

            // manager 6, lane 11, stream 1      
            input   wire                                        std__mgr6__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane11_strm1_data        ,
            output  wire                                        mgr6__std__lane11_strm1_data_valid  ,

            // manager 6, lane 12, stream 0      
            input   wire                                        std__mgr6__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane12_strm0_data        ,
            output  wire                                        mgr6__std__lane12_strm0_data_valid  ,

            // manager 6, lane 12, stream 1      
            input   wire                                        std__mgr6__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane12_strm1_data        ,
            output  wire                                        mgr6__std__lane12_strm1_data_valid  ,

            // manager 6, lane 13, stream 0      
            input   wire                                        std__mgr6__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane13_strm0_data        ,
            output  wire                                        mgr6__std__lane13_strm0_data_valid  ,

            // manager 6, lane 13, stream 1      
            input   wire                                        std__mgr6__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane13_strm1_data        ,
            output  wire                                        mgr6__std__lane13_strm1_data_valid  ,

            // manager 6, lane 14, stream 0      
            input   wire                                        std__mgr6__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane14_strm0_data        ,
            output  wire                                        mgr6__std__lane14_strm0_data_valid  ,

            // manager 6, lane 14, stream 1      
            input   wire                                        std__mgr6__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane14_strm1_data        ,
            output  wire                                        mgr6__std__lane14_strm1_data_valid  ,

            // manager 6, lane 15, stream 0      
            input   wire                                        std__mgr6__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane15_strm0_data        ,
            output  wire                                        mgr6__std__lane15_strm0_data_valid  ,

            // manager 6, lane 15, stream 1      
            input   wire                                        std__mgr6__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane15_strm1_data        ,
            output  wire                                        mgr6__std__lane15_strm1_data_valid  ,

            // manager 6, lane 16, stream 0      
            input   wire                                        std__mgr6__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane16_strm0_data        ,
            output  wire                                        mgr6__std__lane16_strm0_data_valid  ,

            // manager 6, lane 16, stream 1      
            input   wire                                        std__mgr6__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane16_strm1_data        ,
            output  wire                                        mgr6__std__lane16_strm1_data_valid  ,

            // manager 6, lane 17, stream 0      
            input   wire                                        std__mgr6__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane17_strm0_data        ,
            output  wire                                        mgr6__std__lane17_strm0_data_valid  ,

            // manager 6, lane 17, stream 1      
            input   wire                                        std__mgr6__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane17_strm1_data        ,
            output  wire                                        mgr6__std__lane17_strm1_data_valid  ,

            // manager 6, lane 18, stream 0      
            input   wire                                        std__mgr6__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane18_strm0_data        ,
            output  wire                                        mgr6__std__lane18_strm0_data_valid  ,

            // manager 6, lane 18, stream 1      
            input   wire                                        std__mgr6__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane18_strm1_data        ,
            output  wire                                        mgr6__std__lane18_strm1_data_valid  ,

            // manager 6, lane 19, stream 0      
            input   wire                                        std__mgr6__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane19_strm0_data        ,
            output  wire                                        mgr6__std__lane19_strm0_data_valid  ,

            // manager 6, lane 19, stream 1      
            input   wire                                        std__mgr6__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane19_strm1_data        ,
            output  wire                                        mgr6__std__lane19_strm1_data_valid  ,

            // manager 6, lane 20, stream 0      
            input   wire                                        std__mgr6__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane20_strm0_data        ,
            output  wire                                        mgr6__std__lane20_strm0_data_valid  ,

            // manager 6, lane 20, stream 1      
            input   wire                                        std__mgr6__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane20_strm1_data        ,
            output  wire                                        mgr6__std__lane20_strm1_data_valid  ,

            // manager 6, lane 21, stream 0      
            input   wire                                        std__mgr6__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane21_strm0_data        ,
            output  wire                                        mgr6__std__lane21_strm0_data_valid  ,

            // manager 6, lane 21, stream 1      
            input   wire                                        std__mgr6__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane21_strm1_data        ,
            output  wire                                        mgr6__std__lane21_strm1_data_valid  ,

            // manager 6, lane 22, stream 0      
            input   wire                                        std__mgr6__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane22_strm0_data        ,
            output  wire                                        mgr6__std__lane22_strm0_data_valid  ,

            // manager 6, lane 22, stream 1      
            input   wire                                        std__mgr6__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane22_strm1_data        ,
            output  wire                                        mgr6__std__lane22_strm1_data_valid  ,

            // manager 6, lane 23, stream 0      
            input   wire                                        std__mgr6__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane23_strm0_data        ,
            output  wire                                        mgr6__std__lane23_strm0_data_valid  ,

            // manager 6, lane 23, stream 1      
            input   wire                                        std__mgr6__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane23_strm1_data        ,
            output  wire                                        mgr6__std__lane23_strm1_data_valid  ,

            // manager 6, lane 24, stream 0      
            input   wire                                        std__mgr6__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane24_strm0_data        ,
            output  wire                                        mgr6__std__lane24_strm0_data_valid  ,

            // manager 6, lane 24, stream 1      
            input   wire                                        std__mgr6__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane24_strm1_data        ,
            output  wire                                        mgr6__std__lane24_strm1_data_valid  ,

            // manager 6, lane 25, stream 0      
            input   wire                                        std__mgr6__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane25_strm0_data        ,
            output  wire                                        mgr6__std__lane25_strm0_data_valid  ,

            // manager 6, lane 25, stream 1      
            input   wire                                        std__mgr6__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane25_strm1_data        ,
            output  wire                                        mgr6__std__lane25_strm1_data_valid  ,

            // manager 6, lane 26, stream 0      
            input   wire                                        std__mgr6__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane26_strm0_data        ,
            output  wire                                        mgr6__std__lane26_strm0_data_valid  ,

            // manager 6, lane 26, stream 1      
            input   wire                                        std__mgr6__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane26_strm1_data        ,
            output  wire                                        mgr6__std__lane26_strm1_data_valid  ,

            // manager 6, lane 27, stream 0      
            input   wire                                        std__mgr6__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane27_strm0_data        ,
            output  wire                                        mgr6__std__lane27_strm0_data_valid  ,

            // manager 6, lane 27, stream 1      
            input   wire                                        std__mgr6__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane27_strm1_data        ,
            output  wire                                        mgr6__std__lane27_strm1_data_valid  ,

            // manager 6, lane 28, stream 0      
            input   wire                                        std__mgr6__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane28_strm0_data        ,
            output  wire                                        mgr6__std__lane28_strm0_data_valid  ,

            // manager 6, lane 28, stream 1      
            input   wire                                        std__mgr6__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane28_strm1_data        ,
            output  wire                                        mgr6__std__lane28_strm1_data_valid  ,

            // manager 6, lane 29, stream 0      
            input   wire                                        std__mgr6__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane29_strm0_data        ,
            output  wire                                        mgr6__std__lane29_strm0_data_valid  ,

            // manager 6, lane 29, stream 1      
            input   wire                                        std__mgr6__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane29_strm1_data        ,
            output  wire                                        mgr6__std__lane29_strm1_data_valid  ,

            // manager 6, lane 30, stream 0      
            input   wire                                        std__mgr6__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane30_strm0_data        ,
            output  wire                                        mgr6__std__lane30_strm0_data_valid  ,

            // manager 6, lane 30, stream 1      
            input   wire                                        std__mgr6__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane30_strm1_data        ,
            output  wire                                        mgr6__std__lane30_strm1_data_valid  ,

            // manager 6, lane 31, stream 0      
            input   wire                                        std__mgr6__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane31_strm0_data        ,
            output  wire                                        mgr6__std__lane31_strm0_data_valid  ,

            // manager 6, lane 31, stream 1      
            input   wire                                        std__mgr6__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr6__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr6__std__lane31_strm1_data        ,
            output  wire                                        mgr6__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 7, lane 0, stream 0      
            input   wire                                        std__mgr7__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane0_strm0_data        ,
            output  wire                                        mgr7__std__lane0_strm0_data_valid  ,

            // manager 7, lane 0, stream 1      
            input   wire                                        std__mgr7__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane0_strm1_data        ,
            output  wire                                        mgr7__std__lane0_strm1_data_valid  ,

            // manager 7, lane 1, stream 0      
            input   wire                                        std__mgr7__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane1_strm0_data        ,
            output  wire                                        mgr7__std__lane1_strm0_data_valid  ,

            // manager 7, lane 1, stream 1      
            input   wire                                        std__mgr7__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane1_strm1_data        ,
            output  wire                                        mgr7__std__lane1_strm1_data_valid  ,

            // manager 7, lane 2, stream 0      
            input   wire                                        std__mgr7__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane2_strm0_data        ,
            output  wire                                        mgr7__std__lane2_strm0_data_valid  ,

            // manager 7, lane 2, stream 1      
            input   wire                                        std__mgr7__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane2_strm1_data        ,
            output  wire                                        mgr7__std__lane2_strm1_data_valid  ,

            // manager 7, lane 3, stream 0      
            input   wire                                        std__mgr7__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane3_strm0_data        ,
            output  wire                                        mgr7__std__lane3_strm0_data_valid  ,

            // manager 7, lane 3, stream 1      
            input   wire                                        std__mgr7__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane3_strm1_data        ,
            output  wire                                        mgr7__std__lane3_strm1_data_valid  ,

            // manager 7, lane 4, stream 0      
            input   wire                                        std__mgr7__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane4_strm0_data        ,
            output  wire                                        mgr7__std__lane4_strm0_data_valid  ,

            // manager 7, lane 4, stream 1      
            input   wire                                        std__mgr7__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane4_strm1_data        ,
            output  wire                                        mgr7__std__lane4_strm1_data_valid  ,

            // manager 7, lane 5, stream 0      
            input   wire                                        std__mgr7__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane5_strm0_data        ,
            output  wire                                        mgr7__std__lane5_strm0_data_valid  ,

            // manager 7, lane 5, stream 1      
            input   wire                                        std__mgr7__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane5_strm1_data        ,
            output  wire                                        mgr7__std__lane5_strm1_data_valid  ,

            // manager 7, lane 6, stream 0      
            input   wire                                        std__mgr7__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane6_strm0_data        ,
            output  wire                                        mgr7__std__lane6_strm0_data_valid  ,

            // manager 7, lane 6, stream 1      
            input   wire                                        std__mgr7__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane6_strm1_data        ,
            output  wire                                        mgr7__std__lane6_strm1_data_valid  ,

            // manager 7, lane 7, stream 0      
            input   wire                                        std__mgr7__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane7_strm0_data        ,
            output  wire                                        mgr7__std__lane7_strm0_data_valid  ,

            // manager 7, lane 7, stream 1      
            input   wire                                        std__mgr7__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane7_strm1_data        ,
            output  wire                                        mgr7__std__lane7_strm1_data_valid  ,

            // manager 7, lane 8, stream 0      
            input   wire                                        std__mgr7__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane8_strm0_data        ,
            output  wire                                        mgr7__std__lane8_strm0_data_valid  ,

            // manager 7, lane 8, stream 1      
            input   wire                                        std__mgr7__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane8_strm1_data        ,
            output  wire                                        mgr7__std__lane8_strm1_data_valid  ,

            // manager 7, lane 9, stream 0      
            input   wire                                        std__mgr7__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane9_strm0_data        ,
            output  wire                                        mgr7__std__lane9_strm0_data_valid  ,

            // manager 7, lane 9, stream 1      
            input   wire                                        std__mgr7__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane9_strm1_data        ,
            output  wire                                        mgr7__std__lane9_strm1_data_valid  ,

            // manager 7, lane 10, stream 0      
            input   wire                                        std__mgr7__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane10_strm0_data        ,
            output  wire                                        mgr7__std__lane10_strm0_data_valid  ,

            // manager 7, lane 10, stream 1      
            input   wire                                        std__mgr7__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane10_strm1_data        ,
            output  wire                                        mgr7__std__lane10_strm1_data_valid  ,

            // manager 7, lane 11, stream 0      
            input   wire                                        std__mgr7__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane11_strm0_data        ,
            output  wire                                        mgr7__std__lane11_strm0_data_valid  ,

            // manager 7, lane 11, stream 1      
            input   wire                                        std__mgr7__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane11_strm1_data        ,
            output  wire                                        mgr7__std__lane11_strm1_data_valid  ,

            // manager 7, lane 12, stream 0      
            input   wire                                        std__mgr7__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane12_strm0_data        ,
            output  wire                                        mgr7__std__lane12_strm0_data_valid  ,

            // manager 7, lane 12, stream 1      
            input   wire                                        std__mgr7__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane12_strm1_data        ,
            output  wire                                        mgr7__std__lane12_strm1_data_valid  ,

            // manager 7, lane 13, stream 0      
            input   wire                                        std__mgr7__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane13_strm0_data        ,
            output  wire                                        mgr7__std__lane13_strm0_data_valid  ,

            // manager 7, lane 13, stream 1      
            input   wire                                        std__mgr7__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane13_strm1_data        ,
            output  wire                                        mgr7__std__lane13_strm1_data_valid  ,

            // manager 7, lane 14, stream 0      
            input   wire                                        std__mgr7__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane14_strm0_data        ,
            output  wire                                        mgr7__std__lane14_strm0_data_valid  ,

            // manager 7, lane 14, stream 1      
            input   wire                                        std__mgr7__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane14_strm1_data        ,
            output  wire                                        mgr7__std__lane14_strm1_data_valid  ,

            // manager 7, lane 15, stream 0      
            input   wire                                        std__mgr7__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane15_strm0_data        ,
            output  wire                                        mgr7__std__lane15_strm0_data_valid  ,

            // manager 7, lane 15, stream 1      
            input   wire                                        std__mgr7__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane15_strm1_data        ,
            output  wire                                        mgr7__std__lane15_strm1_data_valid  ,

            // manager 7, lane 16, stream 0      
            input   wire                                        std__mgr7__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane16_strm0_data        ,
            output  wire                                        mgr7__std__lane16_strm0_data_valid  ,

            // manager 7, lane 16, stream 1      
            input   wire                                        std__mgr7__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane16_strm1_data        ,
            output  wire                                        mgr7__std__lane16_strm1_data_valid  ,

            // manager 7, lane 17, stream 0      
            input   wire                                        std__mgr7__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane17_strm0_data        ,
            output  wire                                        mgr7__std__lane17_strm0_data_valid  ,

            // manager 7, lane 17, stream 1      
            input   wire                                        std__mgr7__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane17_strm1_data        ,
            output  wire                                        mgr7__std__lane17_strm1_data_valid  ,

            // manager 7, lane 18, stream 0      
            input   wire                                        std__mgr7__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane18_strm0_data        ,
            output  wire                                        mgr7__std__lane18_strm0_data_valid  ,

            // manager 7, lane 18, stream 1      
            input   wire                                        std__mgr7__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane18_strm1_data        ,
            output  wire                                        mgr7__std__lane18_strm1_data_valid  ,

            // manager 7, lane 19, stream 0      
            input   wire                                        std__mgr7__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane19_strm0_data        ,
            output  wire                                        mgr7__std__lane19_strm0_data_valid  ,

            // manager 7, lane 19, stream 1      
            input   wire                                        std__mgr7__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane19_strm1_data        ,
            output  wire                                        mgr7__std__lane19_strm1_data_valid  ,

            // manager 7, lane 20, stream 0      
            input   wire                                        std__mgr7__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane20_strm0_data        ,
            output  wire                                        mgr7__std__lane20_strm0_data_valid  ,

            // manager 7, lane 20, stream 1      
            input   wire                                        std__mgr7__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane20_strm1_data        ,
            output  wire                                        mgr7__std__lane20_strm1_data_valid  ,

            // manager 7, lane 21, stream 0      
            input   wire                                        std__mgr7__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane21_strm0_data        ,
            output  wire                                        mgr7__std__lane21_strm0_data_valid  ,

            // manager 7, lane 21, stream 1      
            input   wire                                        std__mgr7__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane21_strm1_data        ,
            output  wire                                        mgr7__std__lane21_strm1_data_valid  ,

            // manager 7, lane 22, stream 0      
            input   wire                                        std__mgr7__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane22_strm0_data        ,
            output  wire                                        mgr7__std__lane22_strm0_data_valid  ,

            // manager 7, lane 22, stream 1      
            input   wire                                        std__mgr7__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane22_strm1_data        ,
            output  wire                                        mgr7__std__lane22_strm1_data_valid  ,

            // manager 7, lane 23, stream 0      
            input   wire                                        std__mgr7__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane23_strm0_data        ,
            output  wire                                        mgr7__std__lane23_strm0_data_valid  ,

            // manager 7, lane 23, stream 1      
            input   wire                                        std__mgr7__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane23_strm1_data        ,
            output  wire                                        mgr7__std__lane23_strm1_data_valid  ,

            // manager 7, lane 24, stream 0      
            input   wire                                        std__mgr7__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane24_strm0_data        ,
            output  wire                                        mgr7__std__lane24_strm0_data_valid  ,

            // manager 7, lane 24, stream 1      
            input   wire                                        std__mgr7__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane24_strm1_data        ,
            output  wire                                        mgr7__std__lane24_strm1_data_valid  ,

            // manager 7, lane 25, stream 0      
            input   wire                                        std__mgr7__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane25_strm0_data        ,
            output  wire                                        mgr7__std__lane25_strm0_data_valid  ,

            // manager 7, lane 25, stream 1      
            input   wire                                        std__mgr7__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane25_strm1_data        ,
            output  wire                                        mgr7__std__lane25_strm1_data_valid  ,

            // manager 7, lane 26, stream 0      
            input   wire                                        std__mgr7__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane26_strm0_data        ,
            output  wire                                        mgr7__std__lane26_strm0_data_valid  ,

            // manager 7, lane 26, stream 1      
            input   wire                                        std__mgr7__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane26_strm1_data        ,
            output  wire                                        mgr7__std__lane26_strm1_data_valid  ,

            // manager 7, lane 27, stream 0      
            input   wire                                        std__mgr7__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane27_strm0_data        ,
            output  wire                                        mgr7__std__lane27_strm0_data_valid  ,

            // manager 7, lane 27, stream 1      
            input   wire                                        std__mgr7__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane27_strm1_data        ,
            output  wire                                        mgr7__std__lane27_strm1_data_valid  ,

            // manager 7, lane 28, stream 0      
            input   wire                                        std__mgr7__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane28_strm0_data        ,
            output  wire                                        mgr7__std__lane28_strm0_data_valid  ,

            // manager 7, lane 28, stream 1      
            input   wire                                        std__mgr7__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane28_strm1_data        ,
            output  wire                                        mgr7__std__lane28_strm1_data_valid  ,

            // manager 7, lane 29, stream 0      
            input   wire                                        std__mgr7__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane29_strm0_data        ,
            output  wire                                        mgr7__std__lane29_strm0_data_valid  ,

            // manager 7, lane 29, stream 1      
            input   wire                                        std__mgr7__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane29_strm1_data        ,
            output  wire                                        mgr7__std__lane29_strm1_data_valid  ,

            // manager 7, lane 30, stream 0      
            input   wire                                        std__mgr7__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane30_strm0_data        ,
            output  wire                                        mgr7__std__lane30_strm0_data_valid  ,

            // manager 7, lane 30, stream 1      
            input   wire                                        std__mgr7__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane30_strm1_data        ,
            output  wire                                        mgr7__std__lane30_strm1_data_valid  ,

            // manager 7, lane 31, stream 0      
            input   wire                                        std__mgr7__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane31_strm0_data        ,
            output  wire                                        mgr7__std__lane31_strm0_data_valid  ,

            // manager 7, lane 31, stream 1      
            input   wire                                        std__mgr7__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr7__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr7__std__lane31_strm1_data        ,
            output  wire                                        mgr7__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 8, lane 0, stream 0      
            input   wire                                        std__mgr8__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane0_strm0_data        ,
            output  wire                                        mgr8__std__lane0_strm0_data_valid  ,

            // manager 8, lane 0, stream 1      
            input   wire                                        std__mgr8__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane0_strm1_data        ,
            output  wire                                        mgr8__std__lane0_strm1_data_valid  ,

            // manager 8, lane 1, stream 0      
            input   wire                                        std__mgr8__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane1_strm0_data        ,
            output  wire                                        mgr8__std__lane1_strm0_data_valid  ,

            // manager 8, lane 1, stream 1      
            input   wire                                        std__mgr8__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane1_strm1_data        ,
            output  wire                                        mgr8__std__lane1_strm1_data_valid  ,

            // manager 8, lane 2, stream 0      
            input   wire                                        std__mgr8__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane2_strm0_data        ,
            output  wire                                        mgr8__std__lane2_strm0_data_valid  ,

            // manager 8, lane 2, stream 1      
            input   wire                                        std__mgr8__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane2_strm1_data        ,
            output  wire                                        mgr8__std__lane2_strm1_data_valid  ,

            // manager 8, lane 3, stream 0      
            input   wire                                        std__mgr8__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane3_strm0_data        ,
            output  wire                                        mgr8__std__lane3_strm0_data_valid  ,

            // manager 8, lane 3, stream 1      
            input   wire                                        std__mgr8__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane3_strm1_data        ,
            output  wire                                        mgr8__std__lane3_strm1_data_valid  ,

            // manager 8, lane 4, stream 0      
            input   wire                                        std__mgr8__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane4_strm0_data        ,
            output  wire                                        mgr8__std__lane4_strm0_data_valid  ,

            // manager 8, lane 4, stream 1      
            input   wire                                        std__mgr8__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane4_strm1_data        ,
            output  wire                                        mgr8__std__lane4_strm1_data_valid  ,

            // manager 8, lane 5, stream 0      
            input   wire                                        std__mgr8__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane5_strm0_data        ,
            output  wire                                        mgr8__std__lane5_strm0_data_valid  ,

            // manager 8, lane 5, stream 1      
            input   wire                                        std__mgr8__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane5_strm1_data        ,
            output  wire                                        mgr8__std__lane5_strm1_data_valid  ,

            // manager 8, lane 6, stream 0      
            input   wire                                        std__mgr8__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane6_strm0_data        ,
            output  wire                                        mgr8__std__lane6_strm0_data_valid  ,

            // manager 8, lane 6, stream 1      
            input   wire                                        std__mgr8__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane6_strm1_data        ,
            output  wire                                        mgr8__std__lane6_strm1_data_valid  ,

            // manager 8, lane 7, stream 0      
            input   wire                                        std__mgr8__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane7_strm0_data        ,
            output  wire                                        mgr8__std__lane7_strm0_data_valid  ,

            // manager 8, lane 7, stream 1      
            input   wire                                        std__mgr8__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane7_strm1_data        ,
            output  wire                                        mgr8__std__lane7_strm1_data_valid  ,

            // manager 8, lane 8, stream 0      
            input   wire                                        std__mgr8__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane8_strm0_data        ,
            output  wire                                        mgr8__std__lane8_strm0_data_valid  ,

            // manager 8, lane 8, stream 1      
            input   wire                                        std__mgr8__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane8_strm1_data        ,
            output  wire                                        mgr8__std__lane8_strm1_data_valid  ,

            // manager 8, lane 9, stream 0      
            input   wire                                        std__mgr8__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane9_strm0_data        ,
            output  wire                                        mgr8__std__lane9_strm0_data_valid  ,

            // manager 8, lane 9, stream 1      
            input   wire                                        std__mgr8__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane9_strm1_data        ,
            output  wire                                        mgr8__std__lane9_strm1_data_valid  ,

            // manager 8, lane 10, stream 0      
            input   wire                                        std__mgr8__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane10_strm0_data        ,
            output  wire                                        mgr8__std__lane10_strm0_data_valid  ,

            // manager 8, lane 10, stream 1      
            input   wire                                        std__mgr8__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane10_strm1_data        ,
            output  wire                                        mgr8__std__lane10_strm1_data_valid  ,

            // manager 8, lane 11, stream 0      
            input   wire                                        std__mgr8__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane11_strm0_data        ,
            output  wire                                        mgr8__std__lane11_strm0_data_valid  ,

            // manager 8, lane 11, stream 1      
            input   wire                                        std__mgr8__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane11_strm1_data        ,
            output  wire                                        mgr8__std__lane11_strm1_data_valid  ,

            // manager 8, lane 12, stream 0      
            input   wire                                        std__mgr8__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane12_strm0_data        ,
            output  wire                                        mgr8__std__lane12_strm0_data_valid  ,

            // manager 8, lane 12, stream 1      
            input   wire                                        std__mgr8__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane12_strm1_data        ,
            output  wire                                        mgr8__std__lane12_strm1_data_valid  ,

            // manager 8, lane 13, stream 0      
            input   wire                                        std__mgr8__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane13_strm0_data        ,
            output  wire                                        mgr8__std__lane13_strm0_data_valid  ,

            // manager 8, lane 13, stream 1      
            input   wire                                        std__mgr8__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane13_strm1_data        ,
            output  wire                                        mgr8__std__lane13_strm1_data_valid  ,

            // manager 8, lane 14, stream 0      
            input   wire                                        std__mgr8__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane14_strm0_data        ,
            output  wire                                        mgr8__std__lane14_strm0_data_valid  ,

            // manager 8, lane 14, stream 1      
            input   wire                                        std__mgr8__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane14_strm1_data        ,
            output  wire                                        mgr8__std__lane14_strm1_data_valid  ,

            // manager 8, lane 15, stream 0      
            input   wire                                        std__mgr8__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane15_strm0_data        ,
            output  wire                                        mgr8__std__lane15_strm0_data_valid  ,

            // manager 8, lane 15, stream 1      
            input   wire                                        std__mgr8__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane15_strm1_data        ,
            output  wire                                        mgr8__std__lane15_strm1_data_valid  ,

            // manager 8, lane 16, stream 0      
            input   wire                                        std__mgr8__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane16_strm0_data        ,
            output  wire                                        mgr8__std__lane16_strm0_data_valid  ,

            // manager 8, lane 16, stream 1      
            input   wire                                        std__mgr8__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane16_strm1_data        ,
            output  wire                                        mgr8__std__lane16_strm1_data_valid  ,

            // manager 8, lane 17, stream 0      
            input   wire                                        std__mgr8__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane17_strm0_data        ,
            output  wire                                        mgr8__std__lane17_strm0_data_valid  ,

            // manager 8, lane 17, stream 1      
            input   wire                                        std__mgr8__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane17_strm1_data        ,
            output  wire                                        mgr8__std__lane17_strm1_data_valid  ,

            // manager 8, lane 18, stream 0      
            input   wire                                        std__mgr8__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane18_strm0_data        ,
            output  wire                                        mgr8__std__lane18_strm0_data_valid  ,

            // manager 8, lane 18, stream 1      
            input   wire                                        std__mgr8__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane18_strm1_data        ,
            output  wire                                        mgr8__std__lane18_strm1_data_valid  ,

            // manager 8, lane 19, stream 0      
            input   wire                                        std__mgr8__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane19_strm0_data        ,
            output  wire                                        mgr8__std__lane19_strm0_data_valid  ,

            // manager 8, lane 19, stream 1      
            input   wire                                        std__mgr8__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane19_strm1_data        ,
            output  wire                                        mgr8__std__lane19_strm1_data_valid  ,

            // manager 8, lane 20, stream 0      
            input   wire                                        std__mgr8__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane20_strm0_data        ,
            output  wire                                        mgr8__std__lane20_strm0_data_valid  ,

            // manager 8, lane 20, stream 1      
            input   wire                                        std__mgr8__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane20_strm1_data        ,
            output  wire                                        mgr8__std__lane20_strm1_data_valid  ,

            // manager 8, lane 21, stream 0      
            input   wire                                        std__mgr8__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane21_strm0_data        ,
            output  wire                                        mgr8__std__lane21_strm0_data_valid  ,

            // manager 8, lane 21, stream 1      
            input   wire                                        std__mgr8__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane21_strm1_data        ,
            output  wire                                        mgr8__std__lane21_strm1_data_valid  ,

            // manager 8, lane 22, stream 0      
            input   wire                                        std__mgr8__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane22_strm0_data        ,
            output  wire                                        mgr8__std__lane22_strm0_data_valid  ,

            // manager 8, lane 22, stream 1      
            input   wire                                        std__mgr8__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane22_strm1_data        ,
            output  wire                                        mgr8__std__lane22_strm1_data_valid  ,

            // manager 8, lane 23, stream 0      
            input   wire                                        std__mgr8__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane23_strm0_data        ,
            output  wire                                        mgr8__std__lane23_strm0_data_valid  ,

            // manager 8, lane 23, stream 1      
            input   wire                                        std__mgr8__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane23_strm1_data        ,
            output  wire                                        mgr8__std__lane23_strm1_data_valid  ,

            // manager 8, lane 24, stream 0      
            input   wire                                        std__mgr8__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane24_strm0_data        ,
            output  wire                                        mgr8__std__lane24_strm0_data_valid  ,

            // manager 8, lane 24, stream 1      
            input   wire                                        std__mgr8__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane24_strm1_data        ,
            output  wire                                        mgr8__std__lane24_strm1_data_valid  ,

            // manager 8, lane 25, stream 0      
            input   wire                                        std__mgr8__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane25_strm0_data        ,
            output  wire                                        mgr8__std__lane25_strm0_data_valid  ,

            // manager 8, lane 25, stream 1      
            input   wire                                        std__mgr8__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane25_strm1_data        ,
            output  wire                                        mgr8__std__lane25_strm1_data_valid  ,

            // manager 8, lane 26, stream 0      
            input   wire                                        std__mgr8__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane26_strm0_data        ,
            output  wire                                        mgr8__std__lane26_strm0_data_valid  ,

            // manager 8, lane 26, stream 1      
            input   wire                                        std__mgr8__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane26_strm1_data        ,
            output  wire                                        mgr8__std__lane26_strm1_data_valid  ,

            // manager 8, lane 27, stream 0      
            input   wire                                        std__mgr8__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane27_strm0_data        ,
            output  wire                                        mgr8__std__lane27_strm0_data_valid  ,

            // manager 8, lane 27, stream 1      
            input   wire                                        std__mgr8__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane27_strm1_data        ,
            output  wire                                        mgr8__std__lane27_strm1_data_valid  ,

            // manager 8, lane 28, stream 0      
            input   wire                                        std__mgr8__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane28_strm0_data        ,
            output  wire                                        mgr8__std__lane28_strm0_data_valid  ,

            // manager 8, lane 28, stream 1      
            input   wire                                        std__mgr8__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane28_strm1_data        ,
            output  wire                                        mgr8__std__lane28_strm1_data_valid  ,

            // manager 8, lane 29, stream 0      
            input   wire                                        std__mgr8__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane29_strm0_data        ,
            output  wire                                        mgr8__std__lane29_strm0_data_valid  ,

            // manager 8, lane 29, stream 1      
            input   wire                                        std__mgr8__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane29_strm1_data        ,
            output  wire                                        mgr8__std__lane29_strm1_data_valid  ,

            // manager 8, lane 30, stream 0      
            input   wire                                        std__mgr8__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane30_strm0_data        ,
            output  wire                                        mgr8__std__lane30_strm0_data_valid  ,

            // manager 8, lane 30, stream 1      
            input   wire                                        std__mgr8__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane30_strm1_data        ,
            output  wire                                        mgr8__std__lane30_strm1_data_valid  ,

            // manager 8, lane 31, stream 0      
            input   wire                                        std__mgr8__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane31_strm0_data        ,
            output  wire                                        mgr8__std__lane31_strm0_data_valid  ,

            // manager 8, lane 31, stream 1      
            input   wire                                        std__mgr8__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr8__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr8__std__lane31_strm1_data        ,
            output  wire                                        mgr8__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 9, lane 0, stream 0      
            input   wire                                        std__mgr9__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane0_strm0_data        ,
            output  wire                                        mgr9__std__lane0_strm0_data_valid  ,

            // manager 9, lane 0, stream 1      
            input   wire                                        std__mgr9__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane0_strm1_data        ,
            output  wire                                        mgr9__std__lane0_strm1_data_valid  ,

            // manager 9, lane 1, stream 0      
            input   wire                                        std__mgr9__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane1_strm0_data        ,
            output  wire                                        mgr9__std__lane1_strm0_data_valid  ,

            // manager 9, lane 1, stream 1      
            input   wire                                        std__mgr9__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane1_strm1_data        ,
            output  wire                                        mgr9__std__lane1_strm1_data_valid  ,

            // manager 9, lane 2, stream 0      
            input   wire                                        std__mgr9__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane2_strm0_data        ,
            output  wire                                        mgr9__std__lane2_strm0_data_valid  ,

            // manager 9, lane 2, stream 1      
            input   wire                                        std__mgr9__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane2_strm1_data        ,
            output  wire                                        mgr9__std__lane2_strm1_data_valid  ,

            // manager 9, lane 3, stream 0      
            input   wire                                        std__mgr9__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane3_strm0_data        ,
            output  wire                                        mgr9__std__lane3_strm0_data_valid  ,

            // manager 9, lane 3, stream 1      
            input   wire                                        std__mgr9__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane3_strm1_data        ,
            output  wire                                        mgr9__std__lane3_strm1_data_valid  ,

            // manager 9, lane 4, stream 0      
            input   wire                                        std__mgr9__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane4_strm0_data        ,
            output  wire                                        mgr9__std__lane4_strm0_data_valid  ,

            // manager 9, lane 4, stream 1      
            input   wire                                        std__mgr9__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane4_strm1_data        ,
            output  wire                                        mgr9__std__lane4_strm1_data_valid  ,

            // manager 9, lane 5, stream 0      
            input   wire                                        std__mgr9__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane5_strm0_data        ,
            output  wire                                        mgr9__std__lane5_strm0_data_valid  ,

            // manager 9, lane 5, stream 1      
            input   wire                                        std__mgr9__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane5_strm1_data        ,
            output  wire                                        mgr9__std__lane5_strm1_data_valid  ,

            // manager 9, lane 6, stream 0      
            input   wire                                        std__mgr9__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane6_strm0_data        ,
            output  wire                                        mgr9__std__lane6_strm0_data_valid  ,

            // manager 9, lane 6, stream 1      
            input   wire                                        std__mgr9__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane6_strm1_data        ,
            output  wire                                        mgr9__std__lane6_strm1_data_valid  ,

            // manager 9, lane 7, stream 0      
            input   wire                                        std__mgr9__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane7_strm0_data        ,
            output  wire                                        mgr9__std__lane7_strm0_data_valid  ,

            // manager 9, lane 7, stream 1      
            input   wire                                        std__mgr9__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane7_strm1_data        ,
            output  wire                                        mgr9__std__lane7_strm1_data_valid  ,

            // manager 9, lane 8, stream 0      
            input   wire                                        std__mgr9__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane8_strm0_data        ,
            output  wire                                        mgr9__std__lane8_strm0_data_valid  ,

            // manager 9, lane 8, stream 1      
            input   wire                                        std__mgr9__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane8_strm1_data        ,
            output  wire                                        mgr9__std__lane8_strm1_data_valid  ,

            // manager 9, lane 9, stream 0      
            input   wire                                        std__mgr9__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane9_strm0_data        ,
            output  wire                                        mgr9__std__lane9_strm0_data_valid  ,

            // manager 9, lane 9, stream 1      
            input   wire                                        std__mgr9__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane9_strm1_data        ,
            output  wire                                        mgr9__std__lane9_strm1_data_valid  ,

            // manager 9, lane 10, stream 0      
            input   wire                                        std__mgr9__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane10_strm0_data        ,
            output  wire                                        mgr9__std__lane10_strm0_data_valid  ,

            // manager 9, lane 10, stream 1      
            input   wire                                        std__mgr9__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane10_strm1_data        ,
            output  wire                                        mgr9__std__lane10_strm1_data_valid  ,

            // manager 9, lane 11, stream 0      
            input   wire                                        std__mgr9__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane11_strm0_data        ,
            output  wire                                        mgr9__std__lane11_strm0_data_valid  ,

            // manager 9, lane 11, stream 1      
            input   wire                                        std__mgr9__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane11_strm1_data        ,
            output  wire                                        mgr9__std__lane11_strm1_data_valid  ,

            // manager 9, lane 12, stream 0      
            input   wire                                        std__mgr9__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane12_strm0_data        ,
            output  wire                                        mgr9__std__lane12_strm0_data_valid  ,

            // manager 9, lane 12, stream 1      
            input   wire                                        std__mgr9__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane12_strm1_data        ,
            output  wire                                        mgr9__std__lane12_strm1_data_valid  ,

            // manager 9, lane 13, stream 0      
            input   wire                                        std__mgr9__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane13_strm0_data        ,
            output  wire                                        mgr9__std__lane13_strm0_data_valid  ,

            // manager 9, lane 13, stream 1      
            input   wire                                        std__mgr9__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane13_strm1_data        ,
            output  wire                                        mgr9__std__lane13_strm1_data_valid  ,

            // manager 9, lane 14, stream 0      
            input   wire                                        std__mgr9__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane14_strm0_data        ,
            output  wire                                        mgr9__std__lane14_strm0_data_valid  ,

            // manager 9, lane 14, stream 1      
            input   wire                                        std__mgr9__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane14_strm1_data        ,
            output  wire                                        mgr9__std__lane14_strm1_data_valid  ,

            // manager 9, lane 15, stream 0      
            input   wire                                        std__mgr9__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane15_strm0_data        ,
            output  wire                                        mgr9__std__lane15_strm0_data_valid  ,

            // manager 9, lane 15, stream 1      
            input   wire                                        std__mgr9__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane15_strm1_data        ,
            output  wire                                        mgr9__std__lane15_strm1_data_valid  ,

            // manager 9, lane 16, stream 0      
            input   wire                                        std__mgr9__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane16_strm0_data        ,
            output  wire                                        mgr9__std__lane16_strm0_data_valid  ,

            // manager 9, lane 16, stream 1      
            input   wire                                        std__mgr9__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane16_strm1_data        ,
            output  wire                                        mgr9__std__lane16_strm1_data_valid  ,

            // manager 9, lane 17, stream 0      
            input   wire                                        std__mgr9__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane17_strm0_data        ,
            output  wire                                        mgr9__std__lane17_strm0_data_valid  ,

            // manager 9, lane 17, stream 1      
            input   wire                                        std__mgr9__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane17_strm1_data        ,
            output  wire                                        mgr9__std__lane17_strm1_data_valid  ,

            // manager 9, lane 18, stream 0      
            input   wire                                        std__mgr9__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane18_strm0_data        ,
            output  wire                                        mgr9__std__lane18_strm0_data_valid  ,

            // manager 9, lane 18, stream 1      
            input   wire                                        std__mgr9__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane18_strm1_data        ,
            output  wire                                        mgr9__std__lane18_strm1_data_valid  ,

            // manager 9, lane 19, stream 0      
            input   wire                                        std__mgr9__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane19_strm0_data        ,
            output  wire                                        mgr9__std__lane19_strm0_data_valid  ,

            // manager 9, lane 19, stream 1      
            input   wire                                        std__mgr9__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane19_strm1_data        ,
            output  wire                                        mgr9__std__lane19_strm1_data_valid  ,

            // manager 9, lane 20, stream 0      
            input   wire                                        std__mgr9__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane20_strm0_data        ,
            output  wire                                        mgr9__std__lane20_strm0_data_valid  ,

            // manager 9, lane 20, stream 1      
            input   wire                                        std__mgr9__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane20_strm1_data        ,
            output  wire                                        mgr9__std__lane20_strm1_data_valid  ,

            // manager 9, lane 21, stream 0      
            input   wire                                        std__mgr9__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane21_strm0_data        ,
            output  wire                                        mgr9__std__lane21_strm0_data_valid  ,

            // manager 9, lane 21, stream 1      
            input   wire                                        std__mgr9__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane21_strm1_data        ,
            output  wire                                        mgr9__std__lane21_strm1_data_valid  ,

            // manager 9, lane 22, stream 0      
            input   wire                                        std__mgr9__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane22_strm0_data        ,
            output  wire                                        mgr9__std__lane22_strm0_data_valid  ,

            // manager 9, lane 22, stream 1      
            input   wire                                        std__mgr9__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane22_strm1_data        ,
            output  wire                                        mgr9__std__lane22_strm1_data_valid  ,

            // manager 9, lane 23, stream 0      
            input   wire                                        std__mgr9__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane23_strm0_data        ,
            output  wire                                        mgr9__std__lane23_strm0_data_valid  ,

            // manager 9, lane 23, stream 1      
            input   wire                                        std__mgr9__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane23_strm1_data        ,
            output  wire                                        mgr9__std__lane23_strm1_data_valid  ,

            // manager 9, lane 24, stream 0      
            input   wire                                        std__mgr9__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane24_strm0_data        ,
            output  wire                                        mgr9__std__lane24_strm0_data_valid  ,

            // manager 9, lane 24, stream 1      
            input   wire                                        std__mgr9__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane24_strm1_data        ,
            output  wire                                        mgr9__std__lane24_strm1_data_valid  ,

            // manager 9, lane 25, stream 0      
            input   wire                                        std__mgr9__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane25_strm0_data        ,
            output  wire                                        mgr9__std__lane25_strm0_data_valid  ,

            // manager 9, lane 25, stream 1      
            input   wire                                        std__mgr9__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane25_strm1_data        ,
            output  wire                                        mgr9__std__lane25_strm1_data_valid  ,

            // manager 9, lane 26, stream 0      
            input   wire                                        std__mgr9__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane26_strm0_data        ,
            output  wire                                        mgr9__std__lane26_strm0_data_valid  ,

            // manager 9, lane 26, stream 1      
            input   wire                                        std__mgr9__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane26_strm1_data        ,
            output  wire                                        mgr9__std__lane26_strm1_data_valid  ,

            // manager 9, lane 27, stream 0      
            input   wire                                        std__mgr9__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane27_strm0_data        ,
            output  wire                                        mgr9__std__lane27_strm0_data_valid  ,

            // manager 9, lane 27, stream 1      
            input   wire                                        std__mgr9__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane27_strm1_data        ,
            output  wire                                        mgr9__std__lane27_strm1_data_valid  ,

            // manager 9, lane 28, stream 0      
            input   wire                                        std__mgr9__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane28_strm0_data        ,
            output  wire                                        mgr9__std__lane28_strm0_data_valid  ,

            // manager 9, lane 28, stream 1      
            input   wire                                        std__mgr9__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane28_strm1_data        ,
            output  wire                                        mgr9__std__lane28_strm1_data_valid  ,

            // manager 9, lane 29, stream 0      
            input   wire                                        std__mgr9__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane29_strm0_data        ,
            output  wire                                        mgr9__std__lane29_strm0_data_valid  ,

            // manager 9, lane 29, stream 1      
            input   wire                                        std__mgr9__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane29_strm1_data        ,
            output  wire                                        mgr9__std__lane29_strm1_data_valid  ,

            // manager 9, lane 30, stream 0      
            input   wire                                        std__mgr9__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane30_strm0_data        ,
            output  wire                                        mgr9__std__lane30_strm0_data_valid  ,

            // manager 9, lane 30, stream 1      
            input   wire                                        std__mgr9__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane30_strm1_data        ,
            output  wire                                        mgr9__std__lane30_strm1_data_valid  ,

            // manager 9, lane 31, stream 0      
            input   wire                                        std__mgr9__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane31_strm0_data        ,
            output  wire                                        mgr9__std__lane31_strm0_data_valid  ,

            // manager 9, lane 31, stream 1      
            input   wire                                        std__mgr9__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr9__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr9__std__lane31_strm1_data        ,
            output  wire                                        mgr9__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 10, lane 0, stream 0      
            input   wire                                        std__mgr10__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane0_strm0_data        ,
            output  wire                                        mgr10__std__lane0_strm0_data_valid  ,

            // manager 10, lane 0, stream 1      
            input   wire                                        std__mgr10__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane0_strm1_data        ,
            output  wire                                        mgr10__std__lane0_strm1_data_valid  ,

            // manager 10, lane 1, stream 0      
            input   wire                                        std__mgr10__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane1_strm0_data        ,
            output  wire                                        mgr10__std__lane1_strm0_data_valid  ,

            // manager 10, lane 1, stream 1      
            input   wire                                        std__mgr10__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane1_strm1_data        ,
            output  wire                                        mgr10__std__lane1_strm1_data_valid  ,

            // manager 10, lane 2, stream 0      
            input   wire                                        std__mgr10__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane2_strm0_data        ,
            output  wire                                        mgr10__std__lane2_strm0_data_valid  ,

            // manager 10, lane 2, stream 1      
            input   wire                                        std__mgr10__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane2_strm1_data        ,
            output  wire                                        mgr10__std__lane2_strm1_data_valid  ,

            // manager 10, lane 3, stream 0      
            input   wire                                        std__mgr10__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane3_strm0_data        ,
            output  wire                                        mgr10__std__lane3_strm0_data_valid  ,

            // manager 10, lane 3, stream 1      
            input   wire                                        std__mgr10__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane3_strm1_data        ,
            output  wire                                        mgr10__std__lane3_strm1_data_valid  ,

            // manager 10, lane 4, stream 0      
            input   wire                                        std__mgr10__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane4_strm0_data        ,
            output  wire                                        mgr10__std__lane4_strm0_data_valid  ,

            // manager 10, lane 4, stream 1      
            input   wire                                        std__mgr10__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane4_strm1_data        ,
            output  wire                                        mgr10__std__lane4_strm1_data_valid  ,

            // manager 10, lane 5, stream 0      
            input   wire                                        std__mgr10__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane5_strm0_data        ,
            output  wire                                        mgr10__std__lane5_strm0_data_valid  ,

            // manager 10, lane 5, stream 1      
            input   wire                                        std__mgr10__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane5_strm1_data        ,
            output  wire                                        mgr10__std__lane5_strm1_data_valid  ,

            // manager 10, lane 6, stream 0      
            input   wire                                        std__mgr10__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane6_strm0_data        ,
            output  wire                                        mgr10__std__lane6_strm0_data_valid  ,

            // manager 10, lane 6, stream 1      
            input   wire                                        std__mgr10__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane6_strm1_data        ,
            output  wire                                        mgr10__std__lane6_strm1_data_valid  ,

            // manager 10, lane 7, stream 0      
            input   wire                                        std__mgr10__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane7_strm0_data        ,
            output  wire                                        mgr10__std__lane7_strm0_data_valid  ,

            // manager 10, lane 7, stream 1      
            input   wire                                        std__mgr10__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane7_strm1_data        ,
            output  wire                                        mgr10__std__lane7_strm1_data_valid  ,

            // manager 10, lane 8, stream 0      
            input   wire                                        std__mgr10__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane8_strm0_data        ,
            output  wire                                        mgr10__std__lane8_strm0_data_valid  ,

            // manager 10, lane 8, stream 1      
            input   wire                                        std__mgr10__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane8_strm1_data        ,
            output  wire                                        mgr10__std__lane8_strm1_data_valid  ,

            // manager 10, lane 9, stream 0      
            input   wire                                        std__mgr10__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane9_strm0_data        ,
            output  wire                                        mgr10__std__lane9_strm0_data_valid  ,

            // manager 10, lane 9, stream 1      
            input   wire                                        std__mgr10__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane9_strm1_data        ,
            output  wire                                        mgr10__std__lane9_strm1_data_valid  ,

            // manager 10, lane 10, stream 0      
            input   wire                                        std__mgr10__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane10_strm0_data        ,
            output  wire                                        mgr10__std__lane10_strm0_data_valid  ,

            // manager 10, lane 10, stream 1      
            input   wire                                        std__mgr10__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane10_strm1_data        ,
            output  wire                                        mgr10__std__lane10_strm1_data_valid  ,

            // manager 10, lane 11, stream 0      
            input   wire                                        std__mgr10__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane11_strm0_data        ,
            output  wire                                        mgr10__std__lane11_strm0_data_valid  ,

            // manager 10, lane 11, stream 1      
            input   wire                                        std__mgr10__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane11_strm1_data        ,
            output  wire                                        mgr10__std__lane11_strm1_data_valid  ,

            // manager 10, lane 12, stream 0      
            input   wire                                        std__mgr10__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane12_strm0_data        ,
            output  wire                                        mgr10__std__lane12_strm0_data_valid  ,

            // manager 10, lane 12, stream 1      
            input   wire                                        std__mgr10__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane12_strm1_data        ,
            output  wire                                        mgr10__std__lane12_strm1_data_valid  ,

            // manager 10, lane 13, stream 0      
            input   wire                                        std__mgr10__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane13_strm0_data        ,
            output  wire                                        mgr10__std__lane13_strm0_data_valid  ,

            // manager 10, lane 13, stream 1      
            input   wire                                        std__mgr10__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane13_strm1_data        ,
            output  wire                                        mgr10__std__lane13_strm1_data_valid  ,

            // manager 10, lane 14, stream 0      
            input   wire                                        std__mgr10__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane14_strm0_data        ,
            output  wire                                        mgr10__std__lane14_strm0_data_valid  ,

            // manager 10, lane 14, stream 1      
            input   wire                                        std__mgr10__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane14_strm1_data        ,
            output  wire                                        mgr10__std__lane14_strm1_data_valid  ,

            // manager 10, lane 15, stream 0      
            input   wire                                        std__mgr10__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane15_strm0_data        ,
            output  wire                                        mgr10__std__lane15_strm0_data_valid  ,

            // manager 10, lane 15, stream 1      
            input   wire                                        std__mgr10__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane15_strm1_data        ,
            output  wire                                        mgr10__std__lane15_strm1_data_valid  ,

            // manager 10, lane 16, stream 0      
            input   wire                                        std__mgr10__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane16_strm0_data        ,
            output  wire                                        mgr10__std__lane16_strm0_data_valid  ,

            // manager 10, lane 16, stream 1      
            input   wire                                        std__mgr10__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane16_strm1_data        ,
            output  wire                                        mgr10__std__lane16_strm1_data_valid  ,

            // manager 10, lane 17, stream 0      
            input   wire                                        std__mgr10__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane17_strm0_data        ,
            output  wire                                        mgr10__std__lane17_strm0_data_valid  ,

            // manager 10, lane 17, stream 1      
            input   wire                                        std__mgr10__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane17_strm1_data        ,
            output  wire                                        mgr10__std__lane17_strm1_data_valid  ,

            // manager 10, lane 18, stream 0      
            input   wire                                        std__mgr10__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane18_strm0_data        ,
            output  wire                                        mgr10__std__lane18_strm0_data_valid  ,

            // manager 10, lane 18, stream 1      
            input   wire                                        std__mgr10__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane18_strm1_data        ,
            output  wire                                        mgr10__std__lane18_strm1_data_valid  ,

            // manager 10, lane 19, stream 0      
            input   wire                                        std__mgr10__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane19_strm0_data        ,
            output  wire                                        mgr10__std__lane19_strm0_data_valid  ,

            // manager 10, lane 19, stream 1      
            input   wire                                        std__mgr10__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane19_strm1_data        ,
            output  wire                                        mgr10__std__lane19_strm1_data_valid  ,

            // manager 10, lane 20, stream 0      
            input   wire                                        std__mgr10__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane20_strm0_data        ,
            output  wire                                        mgr10__std__lane20_strm0_data_valid  ,

            // manager 10, lane 20, stream 1      
            input   wire                                        std__mgr10__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane20_strm1_data        ,
            output  wire                                        mgr10__std__lane20_strm1_data_valid  ,

            // manager 10, lane 21, stream 0      
            input   wire                                        std__mgr10__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane21_strm0_data        ,
            output  wire                                        mgr10__std__lane21_strm0_data_valid  ,

            // manager 10, lane 21, stream 1      
            input   wire                                        std__mgr10__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane21_strm1_data        ,
            output  wire                                        mgr10__std__lane21_strm1_data_valid  ,

            // manager 10, lane 22, stream 0      
            input   wire                                        std__mgr10__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane22_strm0_data        ,
            output  wire                                        mgr10__std__lane22_strm0_data_valid  ,

            // manager 10, lane 22, stream 1      
            input   wire                                        std__mgr10__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane22_strm1_data        ,
            output  wire                                        mgr10__std__lane22_strm1_data_valid  ,

            // manager 10, lane 23, stream 0      
            input   wire                                        std__mgr10__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane23_strm0_data        ,
            output  wire                                        mgr10__std__lane23_strm0_data_valid  ,

            // manager 10, lane 23, stream 1      
            input   wire                                        std__mgr10__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane23_strm1_data        ,
            output  wire                                        mgr10__std__lane23_strm1_data_valid  ,

            // manager 10, lane 24, stream 0      
            input   wire                                        std__mgr10__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane24_strm0_data        ,
            output  wire                                        mgr10__std__lane24_strm0_data_valid  ,

            // manager 10, lane 24, stream 1      
            input   wire                                        std__mgr10__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane24_strm1_data        ,
            output  wire                                        mgr10__std__lane24_strm1_data_valid  ,

            // manager 10, lane 25, stream 0      
            input   wire                                        std__mgr10__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane25_strm0_data        ,
            output  wire                                        mgr10__std__lane25_strm0_data_valid  ,

            // manager 10, lane 25, stream 1      
            input   wire                                        std__mgr10__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane25_strm1_data        ,
            output  wire                                        mgr10__std__lane25_strm1_data_valid  ,

            // manager 10, lane 26, stream 0      
            input   wire                                        std__mgr10__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane26_strm0_data        ,
            output  wire                                        mgr10__std__lane26_strm0_data_valid  ,

            // manager 10, lane 26, stream 1      
            input   wire                                        std__mgr10__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane26_strm1_data        ,
            output  wire                                        mgr10__std__lane26_strm1_data_valid  ,

            // manager 10, lane 27, stream 0      
            input   wire                                        std__mgr10__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane27_strm0_data        ,
            output  wire                                        mgr10__std__lane27_strm0_data_valid  ,

            // manager 10, lane 27, stream 1      
            input   wire                                        std__mgr10__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane27_strm1_data        ,
            output  wire                                        mgr10__std__lane27_strm1_data_valid  ,

            // manager 10, lane 28, stream 0      
            input   wire                                        std__mgr10__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane28_strm0_data        ,
            output  wire                                        mgr10__std__lane28_strm0_data_valid  ,

            // manager 10, lane 28, stream 1      
            input   wire                                        std__mgr10__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane28_strm1_data        ,
            output  wire                                        mgr10__std__lane28_strm1_data_valid  ,

            // manager 10, lane 29, stream 0      
            input   wire                                        std__mgr10__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane29_strm0_data        ,
            output  wire                                        mgr10__std__lane29_strm0_data_valid  ,

            // manager 10, lane 29, stream 1      
            input   wire                                        std__mgr10__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane29_strm1_data        ,
            output  wire                                        mgr10__std__lane29_strm1_data_valid  ,

            // manager 10, lane 30, stream 0      
            input   wire                                        std__mgr10__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane30_strm0_data        ,
            output  wire                                        mgr10__std__lane30_strm0_data_valid  ,

            // manager 10, lane 30, stream 1      
            input   wire                                        std__mgr10__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane30_strm1_data        ,
            output  wire                                        mgr10__std__lane30_strm1_data_valid  ,

            // manager 10, lane 31, stream 0      
            input   wire                                        std__mgr10__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane31_strm0_data        ,
            output  wire                                        mgr10__std__lane31_strm0_data_valid  ,

            // manager 10, lane 31, stream 1      
            input   wire                                        std__mgr10__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr10__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr10__std__lane31_strm1_data        ,
            output  wire                                        mgr10__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 11, lane 0, stream 0      
            input   wire                                        std__mgr11__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane0_strm0_data        ,
            output  wire                                        mgr11__std__lane0_strm0_data_valid  ,

            // manager 11, lane 0, stream 1      
            input   wire                                        std__mgr11__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane0_strm1_data        ,
            output  wire                                        mgr11__std__lane0_strm1_data_valid  ,

            // manager 11, lane 1, stream 0      
            input   wire                                        std__mgr11__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane1_strm0_data        ,
            output  wire                                        mgr11__std__lane1_strm0_data_valid  ,

            // manager 11, lane 1, stream 1      
            input   wire                                        std__mgr11__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane1_strm1_data        ,
            output  wire                                        mgr11__std__lane1_strm1_data_valid  ,

            // manager 11, lane 2, stream 0      
            input   wire                                        std__mgr11__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane2_strm0_data        ,
            output  wire                                        mgr11__std__lane2_strm0_data_valid  ,

            // manager 11, lane 2, stream 1      
            input   wire                                        std__mgr11__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane2_strm1_data        ,
            output  wire                                        mgr11__std__lane2_strm1_data_valid  ,

            // manager 11, lane 3, stream 0      
            input   wire                                        std__mgr11__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane3_strm0_data        ,
            output  wire                                        mgr11__std__lane3_strm0_data_valid  ,

            // manager 11, lane 3, stream 1      
            input   wire                                        std__mgr11__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane3_strm1_data        ,
            output  wire                                        mgr11__std__lane3_strm1_data_valid  ,

            // manager 11, lane 4, stream 0      
            input   wire                                        std__mgr11__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane4_strm0_data        ,
            output  wire                                        mgr11__std__lane4_strm0_data_valid  ,

            // manager 11, lane 4, stream 1      
            input   wire                                        std__mgr11__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane4_strm1_data        ,
            output  wire                                        mgr11__std__lane4_strm1_data_valid  ,

            // manager 11, lane 5, stream 0      
            input   wire                                        std__mgr11__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane5_strm0_data        ,
            output  wire                                        mgr11__std__lane5_strm0_data_valid  ,

            // manager 11, lane 5, stream 1      
            input   wire                                        std__mgr11__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane5_strm1_data        ,
            output  wire                                        mgr11__std__lane5_strm1_data_valid  ,

            // manager 11, lane 6, stream 0      
            input   wire                                        std__mgr11__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane6_strm0_data        ,
            output  wire                                        mgr11__std__lane6_strm0_data_valid  ,

            // manager 11, lane 6, stream 1      
            input   wire                                        std__mgr11__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane6_strm1_data        ,
            output  wire                                        mgr11__std__lane6_strm1_data_valid  ,

            // manager 11, lane 7, stream 0      
            input   wire                                        std__mgr11__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane7_strm0_data        ,
            output  wire                                        mgr11__std__lane7_strm0_data_valid  ,

            // manager 11, lane 7, stream 1      
            input   wire                                        std__mgr11__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane7_strm1_data        ,
            output  wire                                        mgr11__std__lane7_strm1_data_valid  ,

            // manager 11, lane 8, stream 0      
            input   wire                                        std__mgr11__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane8_strm0_data        ,
            output  wire                                        mgr11__std__lane8_strm0_data_valid  ,

            // manager 11, lane 8, stream 1      
            input   wire                                        std__mgr11__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane8_strm1_data        ,
            output  wire                                        mgr11__std__lane8_strm1_data_valid  ,

            // manager 11, lane 9, stream 0      
            input   wire                                        std__mgr11__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane9_strm0_data        ,
            output  wire                                        mgr11__std__lane9_strm0_data_valid  ,

            // manager 11, lane 9, stream 1      
            input   wire                                        std__mgr11__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane9_strm1_data        ,
            output  wire                                        mgr11__std__lane9_strm1_data_valid  ,

            // manager 11, lane 10, stream 0      
            input   wire                                        std__mgr11__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane10_strm0_data        ,
            output  wire                                        mgr11__std__lane10_strm0_data_valid  ,

            // manager 11, lane 10, stream 1      
            input   wire                                        std__mgr11__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane10_strm1_data        ,
            output  wire                                        mgr11__std__lane10_strm1_data_valid  ,

            // manager 11, lane 11, stream 0      
            input   wire                                        std__mgr11__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane11_strm0_data        ,
            output  wire                                        mgr11__std__lane11_strm0_data_valid  ,

            // manager 11, lane 11, stream 1      
            input   wire                                        std__mgr11__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane11_strm1_data        ,
            output  wire                                        mgr11__std__lane11_strm1_data_valid  ,

            // manager 11, lane 12, stream 0      
            input   wire                                        std__mgr11__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane12_strm0_data        ,
            output  wire                                        mgr11__std__lane12_strm0_data_valid  ,

            // manager 11, lane 12, stream 1      
            input   wire                                        std__mgr11__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane12_strm1_data        ,
            output  wire                                        mgr11__std__lane12_strm1_data_valid  ,

            // manager 11, lane 13, stream 0      
            input   wire                                        std__mgr11__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane13_strm0_data        ,
            output  wire                                        mgr11__std__lane13_strm0_data_valid  ,

            // manager 11, lane 13, stream 1      
            input   wire                                        std__mgr11__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane13_strm1_data        ,
            output  wire                                        mgr11__std__lane13_strm1_data_valid  ,

            // manager 11, lane 14, stream 0      
            input   wire                                        std__mgr11__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane14_strm0_data        ,
            output  wire                                        mgr11__std__lane14_strm0_data_valid  ,

            // manager 11, lane 14, stream 1      
            input   wire                                        std__mgr11__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane14_strm1_data        ,
            output  wire                                        mgr11__std__lane14_strm1_data_valid  ,

            // manager 11, lane 15, stream 0      
            input   wire                                        std__mgr11__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane15_strm0_data        ,
            output  wire                                        mgr11__std__lane15_strm0_data_valid  ,

            // manager 11, lane 15, stream 1      
            input   wire                                        std__mgr11__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane15_strm1_data        ,
            output  wire                                        mgr11__std__lane15_strm1_data_valid  ,

            // manager 11, lane 16, stream 0      
            input   wire                                        std__mgr11__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane16_strm0_data        ,
            output  wire                                        mgr11__std__lane16_strm0_data_valid  ,

            // manager 11, lane 16, stream 1      
            input   wire                                        std__mgr11__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane16_strm1_data        ,
            output  wire                                        mgr11__std__lane16_strm1_data_valid  ,

            // manager 11, lane 17, stream 0      
            input   wire                                        std__mgr11__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane17_strm0_data        ,
            output  wire                                        mgr11__std__lane17_strm0_data_valid  ,

            // manager 11, lane 17, stream 1      
            input   wire                                        std__mgr11__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane17_strm1_data        ,
            output  wire                                        mgr11__std__lane17_strm1_data_valid  ,

            // manager 11, lane 18, stream 0      
            input   wire                                        std__mgr11__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane18_strm0_data        ,
            output  wire                                        mgr11__std__lane18_strm0_data_valid  ,

            // manager 11, lane 18, stream 1      
            input   wire                                        std__mgr11__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane18_strm1_data        ,
            output  wire                                        mgr11__std__lane18_strm1_data_valid  ,

            // manager 11, lane 19, stream 0      
            input   wire                                        std__mgr11__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane19_strm0_data        ,
            output  wire                                        mgr11__std__lane19_strm0_data_valid  ,

            // manager 11, lane 19, stream 1      
            input   wire                                        std__mgr11__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane19_strm1_data        ,
            output  wire                                        mgr11__std__lane19_strm1_data_valid  ,

            // manager 11, lane 20, stream 0      
            input   wire                                        std__mgr11__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane20_strm0_data        ,
            output  wire                                        mgr11__std__lane20_strm0_data_valid  ,

            // manager 11, lane 20, stream 1      
            input   wire                                        std__mgr11__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane20_strm1_data        ,
            output  wire                                        mgr11__std__lane20_strm1_data_valid  ,

            // manager 11, lane 21, stream 0      
            input   wire                                        std__mgr11__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane21_strm0_data        ,
            output  wire                                        mgr11__std__lane21_strm0_data_valid  ,

            // manager 11, lane 21, stream 1      
            input   wire                                        std__mgr11__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane21_strm1_data        ,
            output  wire                                        mgr11__std__lane21_strm1_data_valid  ,

            // manager 11, lane 22, stream 0      
            input   wire                                        std__mgr11__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane22_strm0_data        ,
            output  wire                                        mgr11__std__lane22_strm0_data_valid  ,

            // manager 11, lane 22, stream 1      
            input   wire                                        std__mgr11__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane22_strm1_data        ,
            output  wire                                        mgr11__std__lane22_strm1_data_valid  ,

            // manager 11, lane 23, stream 0      
            input   wire                                        std__mgr11__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane23_strm0_data        ,
            output  wire                                        mgr11__std__lane23_strm0_data_valid  ,

            // manager 11, lane 23, stream 1      
            input   wire                                        std__mgr11__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane23_strm1_data        ,
            output  wire                                        mgr11__std__lane23_strm1_data_valid  ,

            // manager 11, lane 24, stream 0      
            input   wire                                        std__mgr11__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane24_strm0_data        ,
            output  wire                                        mgr11__std__lane24_strm0_data_valid  ,

            // manager 11, lane 24, stream 1      
            input   wire                                        std__mgr11__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane24_strm1_data        ,
            output  wire                                        mgr11__std__lane24_strm1_data_valid  ,

            // manager 11, lane 25, stream 0      
            input   wire                                        std__mgr11__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane25_strm0_data        ,
            output  wire                                        mgr11__std__lane25_strm0_data_valid  ,

            // manager 11, lane 25, stream 1      
            input   wire                                        std__mgr11__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane25_strm1_data        ,
            output  wire                                        mgr11__std__lane25_strm1_data_valid  ,

            // manager 11, lane 26, stream 0      
            input   wire                                        std__mgr11__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane26_strm0_data        ,
            output  wire                                        mgr11__std__lane26_strm0_data_valid  ,

            // manager 11, lane 26, stream 1      
            input   wire                                        std__mgr11__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane26_strm1_data        ,
            output  wire                                        mgr11__std__lane26_strm1_data_valid  ,

            // manager 11, lane 27, stream 0      
            input   wire                                        std__mgr11__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane27_strm0_data        ,
            output  wire                                        mgr11__std__lane27_strm0_data_valid  ,

            // manager 11, lane 27, stream 1      
            input   wire                                        std__mgr11__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane27_strm1_data        ,
            output  wire                                        mgr11__std__lane27_strm1_data_valid  ,

            // manager 11, lane 28, stream 0      
            input   wire                                        std__mgr11__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane28_strm0_data        ,
            output  wire                                        mgr11__std__lane28_strm0_data_valid  ,

            // manager 11, lane 28, stream 1      
            input   wire                                        std__mgr11__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane28_strm1_data        ,
            output  wire                                        mgr11__std__lane28_strm1_data_valid  ,

            // manager 11, lane 29, stream 0      
            input   wire                                        std__mgr11__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane29_strm0_data        ,
            output  wire                                        mgr11__std__lane29_strm0_data_valid  ,

            // manager 11, lane 29, stream 1      
            input   wire                                        std__mgr11__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane29_strm1_data        ,
            output  wire                                        mgr11__std__lane29_strm1_data_valid  ,

            // manager 11, lane 30, stream 0      
            input   wire                                        std__mgr11__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane30_strm0_data        ,
            output  wire                                        mgr11__std__lane30_strm0_data_valid  ,

            // manager 11, lane 30, stream 1      
            input   wire                                        std__mgr11__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane30_strm1_data        ,
            output  wire                                        mgr11__std__lane30_strm1_data_valid  ,

            // manager 11, lane 31, stream 0      
            input   wire                                        std__mgr11__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane31_strm0_data        ,
            output  wire                                        mgr11__std__lane31_strm0_data_valid  ,

            // manager 11, lane 31, stream 1      
            input   wire                                        std__mgr11__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr11__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr11__std__lane31_strm1_data        ,
            output  wire                                        mgr11__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 12, lane 0, stream 0      
            input   wire                                        std__mgr12__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane0_strm0_data        ,
            output  wire                                        mgr12__std__lane0_strm0_data_valid  ,

            // manager 12, lane 0, stream 1      
            input   wire                                        std__mgr12__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane0_strm1_data        ,
            output  wire                                        mgr12__std__lane0_strm1_data_valid  ,

            // manager 12, lane 1, stream 0      
            input   wire                                        std__mgr12__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane1_strm0_data        ,
            output  wire                                        mgr12__std__lane1_strm0_data_valid  ,

            // manager 12, lane 1, stream 1      
            input   wire                                        std__mgr12__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane1_strm1_data        ,
            output  wire                                        mgr12__std__lane1_strm1_data_valid  ,

            // manager 12, lane 2, stream 0      
            input   wire                                        std__mgr12__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane2_strm0_data        ,
            output  wire                                        mgr12__std__lane2_strm0_data_valid  ,

            // manager 12, lane 2, stream 1      
            input   wire                                        std__mgr12__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane2_strm1_data        ,
            output  wire                                        mgr12__std__lane2_strm1_data_valid  ,

            // manager 12, lane 3, stream 0      
            input   wire                                        std__mgr12__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane3_strm0_data        ,
            output  wire                                        mgr12__std__lane3_strm0_data_valid  ,

            // manager 12, lane 3, stream 1      
            input   wire                                        std__mgr12__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane3_strm1_data        ,
            output  wire                                        mgr12__std__lane3_strm1_data_valid  ,

            // manager 12, lane 4, stream 0      
            input   wire                                        std__mgr12__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane4_strm0_data        ,
            output  wire                                        mgr12__std__lane4_strm0_data_valid  ,

            // manager 12, lane 4, stream 1      
            input   wire                                        std__mgr12__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane4_strm1_data        ,
            output  wire                                        mgr12__std__lane4_strm1_data_valid  ,

            // manager 12, lane 5, stream 0      
            input   wire                                        std__mgr12__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane5_strm0_data        ,
            output  wire                                        mgr12__std__lane5_strm0_data_valid  ,

            // manager 12, lane 5, stream 1      
            input   wire                                        std__mgr12__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane5_strm1_data        ,
            output  wire                                        mgr12__std__lane5_strm1_data_valid  ,

            // manager 12, lane 6, stream 0      
            input   wire                                        std__mgr12__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane6_strm0_data        ,
            output  wire                                        mgr12__std__lane6_strm0_data_valid  ,

            // manager 12, lane 6, stream 1      
            input   wire                                        std__mgr12__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane6_strm1_data        ,
            output  wire                                        mgr12__std__lane6_strm1_data_valid  ,

            // manager 12, lane 7, stream 0      
            input   wire                                        std__mgr12__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane7_strm0_data        ,
            output  wire                                        mgr12__std__lane7_strm0_data_valid  ,

            // manager 12, lane 7, stream 1      
            input   wire                                        std__mgr12__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane7_strm1_data        ,
            output  wire                                        mgr12__std__lane7_strm1_data_valid  ,

            // manager 12, lane 8, stream 0      
            input   wire                                        std__mgr12__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane8_strm0_data        ,
            output  wire                                        mgr12__std__lane8_strm0_data_valid  ,

            // manager 12, lane 8, stream 1      
            input   wire                                        std__mgr12__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane8_strm1_data        ,
            output  wire                                        mgr12__std__lane8_strm1_data_valid  ,

            // manager 12, lane 9, stream 0      
            input   wire                                        std__mgr12__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane9_strm0_data        ,
            output  wire                                        mgr12__std__lane9_strm0_data_valid  ,

            // manager 12, lane 9, stream 1      
            input   wire                                        std__mgr12__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane9_strm1_data        ,
            output  wire                                        mgr12__std__lane9_strm1_data_valid  ,

            // manager 12, lane 10, stream 0      
            input   wire                                        std__mgr12__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane10_strm0_data        ,
            output  wire                                        mgr12__std__lane10_strm0_data_valid  ,

            // manager 12, lane 10, stream 1      
            input   wire                                        std__mgr12__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane10_strm1_data        ,
            output  wire                                        mgr12__std__lane10_strm1_data_valid  ,

            // manager 12, lane 11, stream 0      
            input   wire                                        std__mgr12__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane11_strm0_data        ,
            output  wire                                        mgr12__std__lane11_strm0_data_valid  ,

            // manager 12, lane 11, stream 1      
            input   wire                                        std__mgr12__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane11_strm1_data        ,
            output  wire                                        mgr12__std__lane11_strm1_data_valid  ,

            // manager 12, lane 12, stream 0      
            input   wire                                        std__mgr12__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane12_strm0_data        ,
            output  wire                                        mgr12__std__lane12_strm0_data_valid  ,

            // manager 12, lane 12, stream 1      
            input   wire                                        std__mgr12__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane12_strm1_data        ,
            output  wire                                        mgr12__std__lane12_strm1_data_valid  ,

            // manager 12, lane 13, stream 0      
            input   wire                                        std__mgr12__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane13_strm0_data        ,
            output  wire                                        mgr12__std__lane13_strm0_data_valid  ,

            // manager 12, lane 13, stream 1      
            input   wire                                        std__mgr12__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane13_strm1_data        ,
            output  wire                                        mgr12__std__lane13_strm1_data_valid  ,

            // manager 12, lane 14, stream 0      
            input   wire                                        std__mgr12__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane14_strm0_data        ,
            output  wire                                        mgr12__std__lane14_strm0_data_valid  ,

            // manager 12, lane 14, stream 1      
            input   wire                                        std__mgr12__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane14_strm1_data        ,
            output  wire                                        mgr12__std__lane14_strm1_data_valid  ,

            // manager 12, lane 15, stream 0      
            input   wire                                        std__mgr12__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane15_strm0_data        ,
            output  wire                                        mgr12__std__lane15_strm0_data_valid  ,

            // manager 12, lane 15, stream 1      
            input   wire                                        std__mgr12__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane15_strm1_data        ,
            output  wire                                        mgr12__std__lane15_strm1_data_valid  ,

            // manager 12, lane 16, stream 0      
            input   wire                                        std__mgr12__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane16_strm0_data        ,
            output  wire                                        mgr12__std__lane16_strm0_data_valid  ,

            // manager 12, lane 16, stream 1      
            input   wire                                        std__mgr12__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane16_strm1_data        ,
            output  wire                                        mgr12__std__lane16_strm1_data_valid  ,

            // manager 12, lane 17, stream 0      
            input   wire                                        std__mgr12__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane17_strm0_data        ,
            output  wire                                        mgr12__std__lane17_strm0_data_valid  ,

            // manager 12, lane 17, stream 1      
            input   wire                                        std__mgr12__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane17_strm1_data        ,
            output  wire                                        mgr12__std__lane17_strm1_data_valid  ,

            // manager 12, lane 18, stream 0      
            input   wire                                        std__mgr12__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane18_strm0_data        ,
            output  wire                                        mgr12__std__lane18_strm0_data_valid  ,

            // manager 12, lane 18, stream 1      
            input   wire                                        std__mgr12__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane18_strm1_data        ,
            output  wire                                        mgr12__std__lane18_strm1_data_valid  ,

            // manager 12, lane 19, stream 0      
            input   wire                                        std__mgr12__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane19_strm0_data        ,
            output  wire                                        mgr12__std__lane19_strm0_data_valid  ,

            // manager 12, lane 19, stream 1      
            input   wire                                        std__mgr12__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane19_strm1_data        ,
            output  wire                                        mgr12__std__lane19_strm1_data_valid  ,

            // manager 12, lane 20, stream 0      
            input   wire                                        std__mgr12__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane20_strm0_data        ,
            output  wire                                        mgr12__std__lane20_strm0_data_valid  ,

            // manager 12, lane 20, stream 1      
            input   wire                                        std__mgr12__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane20_strm1_data        ,
            output  wire                                        mgr12__std__lane20_strm1_data_valid  ,

            // manager 12, lane 21, stream 0      
            input   wire                                        std__mgr12__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane21_strm0_data        ,
            output  wire                                        mgr12__std__lane21_strm0_data_valid  ,

            // manager 12, lane 21, stream 1      
            input   wire                                        std__mgr12__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane21_strm1_data        ,
            output  wire                                        mgr12__std__lane21_strm1_data_valid  ,

            // manager 12, lane 22, stream 0      
            input   wire                                        std__mgr12__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane22_strm0_data        ,
            output  wire                                        mgr12__std__lane22_strm0_data_valid  ,

            // manager 12, lane 22, stream 1      
            input   wire                                        std__mgr12__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane22_strm1_data        ,
            output  wire                                        mgr12__std__lane22_strm1_data_valid  ,

            // manager 12, lane 23, stream 0      
            input   wire                                        std__mgr12__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane23_strm0_data        ,
            output  wire                                        mgr12__std__lane23_strm0_data_valid  ,

            // manager 12, lane 23, stream 1      
            input   wire                                        std__mgr12__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane23_strm1_data        ,
            output  wire                                        mgr12__std__lane23_strm1_data_valid  ,

            // manager 12, lane 24, stream 0      
            input   wire                                        std__mgr12__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane24_strm0_data        ,
            output  wire                                        mgr12__std__lane24_strm0_data_valid  ,

            // manager 12, lane 24, stream 1      
            input   wire                                        std__mgr12__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane24_strm1_data        ,
            output  wire                                        mgr12__std__lane24_strm1_data_valid  ,

            // manager 12, lane 25, stream 0      
            input   wire                                        std__mgr12__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane25_strm0_data        ,
            output  wire                                        mgr12__std__lane25_strm0_data_valid  ,

            // manager 12, lane 25, stream 1      
            input   wire                                        std__mgr12__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane25_strm1_data        ,
            output  wire                                        mgr12__std__lane25_strm1_data_valid  ,

            // manager 12, lane 26, stream 0      
            input   wire                                        std__mgr12__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane26_strm0_data        ,
            output  wire                                        mgr12__std__lane26_strm0_data_valid  ,

            // manager 12, lane 26, stream 1      
            input   wire                                        std__mgr12__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane26_strm1_data        ,
            output  wire                                        mgr12__std__lane26_strm1_data_valid  ,

            // manager 12, lane 27, stream 0      
            input   wire                                        std__mgr12__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane27_strm0_data        ,
            output  wire                                        mgr12__std__lane27_strm0_data_valid  ,

            // manager 12, lane 27, stream 1      
            input   wire                                        std__mgr12__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane27_strm1_data        ,
            output  wire                                        mgr12__std__lane27_strm1_data_valid  ,

            // manager 12, lane 28, stream 0      
            input   wire                                        std__mgr12__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane28_strm0_data        ,
            output  wire                                        mgr12__std__lane28_strm0_data_valid  ,

            // manager 12, lane 28, stream 1      
            input   wire                                        std__mgr12__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane28_strm1_data        ,
            output  wire                                        mgr12__std__lane28_strm1_data_valid  ,

            // manager 12, lane 29, stream 0      
            input   wire                                        std__mgr12__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane29_strm0_data        ,
            output  wire                                        mgr12__std__lane29_strm0_data_valid  ,

            // manager 12, lane 29, stream 1      
            input   wire                                        std__mgr12__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane29_strm1_data        ,
            output  wire                                        mgr12__std__lane29_strm1_data_valid  ,

            // manager 12, lane 30, stream 0      
            input   wire                                        std__mgr12__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane30_strm0_data        ,
            output  wire                                        mgr12__std__lane30_strm0_data_valid  ,

            // manager 12, lane 30, stream 1      
            input   wire                                        std__mgr12__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane30_strm1_data        ,
            output  wire                                        mgr12__std__lane30_strm1_data_valid  ,

            // manager 12, lane 31, stream 0      
            input   wire                                        std__mgr12__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane31_strm0_data        ,
            output  wire                                        mgr12__std__lane31_strm0_data_valid  ,

            // manager 12, lane 31, stream 1      
            input   wire                                        std__mgr12__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr12__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr12__std__lane31_strm1_data        ,
            output  wire                                        mgr12__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 13, lane 0, stream 0      
            input   wire                                        std__mgr13__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane0_strm0_data        ,
            output  wire                                        mgr13__std__lane0_strm0_data_valid  ,

            // manager 13, lane 0, stream 1      
            input   wire                                        std__mgr13__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane0_strm1_data        ,
            output  wire                                        mgr13__std__lane0_strm1_data_valid  ,

            // manager 13, lane 1, stream 0      
            input   wire                                        std__mgr13__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane1_strm0_data        ,
            output  wire                                        mgr13__std__lane1_strm0_data_valid  ,

            // manager 13, lane 1, stream 1      
            input   wire                                        std__mgr13__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane1_strm1_data        ,
            output  wire                                        mgr13__std__lane1_strm1_data_valid  ,

            // manager 13, lane 2, stream 0      
            input   wire                                        std__mgr13__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane2_strm0_data        ,
            output  wire                                        mgr13__std__lane2_strm0_data_valid  ,

            // manager 13, lane 2, stream 1      
            input   wire                                        std__mgr13__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane2_strm1_data        ,
            output  wire                                        mgr13__std__lane2_strm1_data_valid  ,

            // manager 13, lane 3, stream 0      
            input   wire                                        std__mgr13__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane3_strm0_data        ,
            output  wire                                        mgr13__std__lane3_strm0_data_valid  ,

            // manager 13, lane 3, stream 1      
            input   wire                                        std__mgr13__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane3_strm1_data        ,
            output  wire                                        mgr13__std__lane3_strm1_data_valid  ,

            // manager 13, lane 4, stream 0      
            input   wire                                        std__mgr13__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane4_strm0_data        ,
            output  wire                                        mgr13__std__lane4_strm0_data_valid  ,

            // manager 13, lane 4, stream 1      
            input   wire                                        std__mgr13__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane4_strm1_data        ,
            output  wire                                        mgr13__std__lane4_strm1_data_valid  ,

            // manager 13, lane 5, stream 0      
            input   wire                                        std__mgr13__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane5_strm0_data        ,
            output  wire                                        mgr13__std__lane5_strm0_data_valid  ,

            // manager 13, lane 5, stream 1      
            input   wire                                        std__mgr13__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane5_strm1_data        ,
            output  wire                                        mgr13__std__lane5_strm1_data_valid  ,

            // manager 13, lane 6, stream 0      
            input   wire                                        std__mgr13__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane6_strm0_data        ,
            output  wire                                        mgr13__std__lane6_strm0_data_valid  ,

            // manager 13, lane 6, stream 1      
            input   wire                                        std__mgr13__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane6_strm1_data        ,
            output  wire                                        mgr13__std__lane6_strm1_data_valid  ,

            // manager 13, lane 7, stream 0      
            input   wire                                        std__mgr13__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane7_strm0_data        ,
            output  wire                                        mgr13__std__lane7_strm0_data_valid  ,

            // manager 13, lane 7, stream 1      
            input   wire                                        std__mgr13__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane7_strm1_data        ,
            output  wire                                        mgr13__std__lane7_strm1_data_valid  ,

            // manager 13, lane 8, stream 0      
            input   wire                                        std__mgr13__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane8_strm0_data        ,
            output  wire                                        mgr13__std__lane8_strm0_data_valid  ,

            // manager 13, lane 8, stream 1      
            input   wire                                        std__mgr13__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane8_strm1_data        ,
            output  wire                                        mgr13__std__lane8_strm1_data_valid  ,

            // manager 13, lane 9, stream 0      
            input   wire                                        std__mgr13__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane9_strm0_data        ,
            output  wire                                        mgr13__std__lane9_strm0_data_valid  ,

            // manager 13, lane 9, stream 1      
            input   wire                                        std__mgr13__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane9_strm1_data        ,
            output  wire                                        mgr13__std__lane9_strm1_data_valid  ,

            // manager 13, lane 10, stream 0      
            input   wire                                        std__mgr13__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane10_strm0_data        ,
            output  wire                                        mgr13__std__lane10_strm0_data_valid  ,

            // manager 13, lane 10, stream 1      
            input   wire                                        std__mgr13__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane10_strm1_data        ,
            output  wire                                        mgr13__std__lane10_strm1_data_valid  ,

            // manager 13, lane 11, stream 0      
            input   wire                                        std__mgr13__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane11_strm0_data        ,
            output  wire                                        mgr13__std__lane11_strm0_data_valid  ,

            // manager 13, lane 11, stream 1      
            input   wire                                        std__mgr13__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane11_strm1_data        ,
            output  wire                                        mgr13__std__lane11_strm1_data_valid  ,

            // manager 13, lane 12, stream 0      
            input   wire                                        std__mgr13__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane12_strm0_data        ,
            output  wire                                        mgr13__std__lane12_strm0_data_valid  ,

            // manager 13, lane 12, stream 1      
            input   wire                                        std__mgr13__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane12_strm1_data        ,
            output  wire                                        mgr13__std__lane12_strm1_data_valid  ,

            // manager 13, lane 13, stream 0      
            input   wire                                        std__mgr13__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane13_strm0_data        ,
            output  wire                                        mgr13__std__lane13_strm0_data_valid  ,

            // manager 13, lane 13, stream 1      
            input   wire                                        std__mgr13__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane13_strm1_data        ,
            output  wire                                        mgr13__std__lane13_strm1_data_valid  ,

            // manager 13, lane 14, stream 0      
            input   wire                                        std__mgr13__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane14_strm0_data        ,
            output  wire                                        mgr13__std__lane14_strm0_data_valid  ,

            // manager 13, lane 14, stream 1      
            input   wire                                        std__mgr13__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane14_strm1_data        ,
            output  wire                                        mgr13__std__lane14_strm1_data_valid  ,

            // manager 13, lane 15, stream 0      
            input   wire                                        std__mgr13__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane15_strm0_data        ,
            output  wire                                        mgr13__std__lane15_strm0_data_valid  ,

            // manager 13, lane 15, stream 1      
            input   wire                                        std__mgr13__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane15_strm1_data        ,
            output  wire                                        mgr13__std__lane15_strm1_data_valid  ,

            // manager 13, lane 16, stream 0      
            input   wire                                        std__mgr13__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane16_strm0_data        ,
            output  wire                                        mgr13__std__lane16_strm0_data_valid  ,

            // manager 13, lane 16, stream 1      
            input   wire                                        std__mgr13__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane16_strm1_data        ,
            output  wire                                        mgr13__std__lane16_strm1_data_valid  ,

            // manager 13, lane 17, stream 0      
            input   wire                                        std__mgr13__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane17_strm0_data        ,
            output  wire                                        mgr13__std__lane17_strm0_data_valid  ,

            // manager 13, lane 17, stream 1      
            input   wire                                        std__mgr13__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane17_strm1_data        ,
            output  wire                                        mgr13__std__lane17_strm1_data_valid  ,

            // manager 13, lane 18, stream 0      
            input   wire                                        std__mgr13__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane18_strm0_data        ,
            output  wire                                        mgr13__std__lane18_strm0_data_valid  ,

            // manager 13, lane 18, stream 1      
            input   wire                                        std__mgr13__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane18_strm1_data        ,
            output  wire                                        mgr13__std__lane18_strm1_data_valid  ,

            // manager 13, lane 19, stream 0      
            input   wire                                        std__mgr13__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane19_strm0_data        ,
            output  wire                                        mgr13__std__lane19_strm0_data_valid  ,

            // manager 13, lane 19, stream 1      
            input   wire                                        std__mgr13__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane19_strm1_data        ,
            output  wire                                        mgr13__std__lane19_strm1_data_valid  ,

            // manager 13, lane 20, stream 0      
            input   wire                                        std__mgr13__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane20_strm0_data        ,
            output  wire                                        mgr13__std__lane20_strm0_data_valid  ,

            // manager 13, lane 20, stream 1      
            input   wire                                        std__mgr13__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane20_strm1_data        ,
            output  wire                                        mgr13__std__lane20_strm1_data_valid  ,

            // manager 13, lane 21, stream 0      
            input   wire                                        std__mgr13__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane21_strm0_data        ,
            output  wire                                        mgr13__std__lane21_strm0_data_valid  ,

            // manager 13, lane 21, stream 1      
            input   wire                                        std__mgr13__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane21_strm1_data        ,
            output  wire                                        mgr13__std__lane21_strm1_data_valid  ,

            // manager 13, lane 22, stream 0      
            input   wire                                        std__mgr13__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane22_strm0_data        ,
            output  wire                                        mgr13__std__lane22_strm0_data_valid  ,

            // manager 13, lane 22, stream 1      
            input   wire                                        std__mgr13__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane22_strm1_data        ,
            output  wire                                        mgr13__std__lane22_strm1_data_valid  ,

            // manager 13, lane 23, stream 0      
            input   wire                                        std__mgr13__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane23_strm0_data        ,
            output  wire                                        mgr13__std__lane23_strm0_data_valid  ,

            // manager 13, lane 23, stream 1      
            input   wire                                        std__mgr13__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane23_strm1_data        ,
            output  wire                                        mgr13__std__lane23_strm1_data_valid  ,

            // manager 13, lane 24, stream 0      
            input   wire                                        std__mgr13__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane24_strm0_data        ,
            output  wire                                        mgr13__std__lane24_strm0_data_valid  ,

            // manager 13, lane 24, stream 1      
            input   wire                                        std__mgr13__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane24_strm1_data        ,
            output  wire                                        mgr13__std__lane24_strm1_data_valid  ,

            // manager 13, lane 25, stream 0      
            input   wire                                        std__mgr13__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane25_strm0_data        ,
            output  wire                                        mgr13__std__lane25_strm0_data_valid  ,

            // manager 13, lane 25, stream 1      
            input   wire                                        std__mgr13__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane25_strm1_data        ,
            output  wire                                        mgr13__std__lane25_strm1_data_valid  ,

            // manager 13, lane 26, stream 0      
            input   wire                                        std__mgr13__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane26_strm0_data        ,
            output  wire                                        mgr13__std__lane26_strm0_data_valid  ,

            // manager 13, lane 26, stream 1      
            input   wire                                        std__mgr13__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane26_strm1_data        ,
            output  wire                                        mgr13__std__lane26_strm1_data_valid  ,

            // manager 13, lane 27, stream 0      
            input   wire                                        std__mgr13__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane27_strm0_data        ,
            output  wire                                        mgr13__std__lane27_strm0_data_valid  ,

            // manager 13, lane 27, stream 1      
            input   wire                                        std__mgr13__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane27_strm1_data        ,
            output  wire                                        mgr13__std__lane27_strm1_data_valid  ,

            // manager 13, lane 28, stream 0      
            input   wire                                        std__mgr13__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane28_strm0_data        ,
            output  wire                                        mgr13__std__lane28_strm0_data_valid  ,

            // manager 13, lane 28, stream 1      
            input   wire                                        std__mgr13__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane28_strm1_data        ,
            output  wire                                        mgr13__std__lane28_strm1_data_valid  ,

            // manager 13, lane 29, stream 0      
            input   wire                                        std__mgr13__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane29_strm0_data        ,
            output  wire                                        mgr13__std__lane29_strm0_data_valid  ,

            // manager 13, lane 29, stream 1      
            input   wire                                        std__mgr13__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane29_strm1_data        ,
            output  wire                                        mgr13__std__lane29_strm1_data_valid  ,

            // manager 13, lane 30, stream 0      
            input   wire                                        std__mgr13__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane30_strm0_data        ,
            output  wire                                        mgr13__std__lane30_strm0_data_valid  ,

            // manager 13, lane 30, stream 1      
            input   wire                                        std__mgr13__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane30_strm1_data        ,
            output  wire                                        mgr13__std__lane30_strm1_data_valid  ,

            // manager 13, lane 31, stream 0      
            input   wire                                        std__mgr13__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane31_strm0_data        ,
            output  wire                                        mgr13__std__lane31_strm0_data_valid  ,

            // manager 13, lane 31, stream 1      
            input   wire                                        std__mgr13__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr13__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr13__std__lane31_strm1_data        ,
            output  wire                                        mgr13__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 14, lane 0, stream 0      
            input   wire                                        std__mgr14__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane0_strm0_data        ,
            output  wire                                        mgr14__std__lane0_strm0_data_valid  ,

            // manager 14, lane 0, stream 1      
            input   wire                                        std__mgr14__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane0_strm1_data        ,
            output  wire                                        mgr14__std__lane0_strm1_data_valid  ,

            // manager 14, lane 1, stream 0      
            input   wire                                        std__mgr14__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane1_strm0_data        ,
            output  wire                                        mgr14__std__lane1_strm0_data_valid  ,

            // manager 14, lane 1, stream 1      
            input   wire                                        std__mgr14__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane1_strm1_data        ,
            output  wire                                        mgr14__std__lane1_strm1_data_valid  ,

            // manager 14, lane 2, stream 0      
            input   wire                                        std__mgr14__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane2_strm0_data        ,
            output  wire                                        mgr14__std__lane2_strm0_data_valid  ,

            // manager 14, lane 2, stream 1      
            input   wire                                        std__mgr14__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane2_strm1_data        ,
            output  wire                                        mgr14__std__lane2_strm1_data_valid  ,

            // manager 14, lane 3, stream 0      
            input   wire                                        std__mgr14__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane3_strm0_data        ,
            output  wire                                        mgr14__std__lane3_strm0_data_valid  ,

            // manager 14, lane 3, stream 1      
            input   wire                                        std__mgr14__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane3_strm1_data        ,
            output  wire                                        mgr14__std__lane3_strm1_data_valid  ,

            // manager 14, lane 4, stream 0      
            input   wire                                        std__mgr14__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane4_strm0_data        ,
            output  wire                                        mgr14__std__lane4_strm0_data_valid  ,

            // manager 14, lane 4, stream 1      
            input   wire                                        std__mgr14__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane4_strm1_data        ,
            output  wire                                        mgr14__std__lane4_strm1_data_valid  ,

            // manager 14, lane 5, stream 0      
            input   wire                                        std__mgr14__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane5_strm0_data        ,
            output  wire                                        mgr14__std__lane5_strm0_data_valid  ,

            // manager 14, lane 5, stream 1      
            input   wire                                        std__mgr14__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane5_strm1_data        ,
            output  wire                                        mgr14__std__lane5_strm1_data_valid  ,

            // manager 14, lane 6, stream 0      
            input   wire                                        std__mgr14__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane6_strm0_data        ,
            output  wire                                        mgr14__std__lane6_strm0_data_valid  ,

            // manager 14, lane 6, stream 1      
            input   wire                                        std__mgr14__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane6_strm1_data        ,
            output  wire                                        mgr14__std__lane6_strm1_data_valid  ,

            // manager 14, lane 7, stream 0      
            input   wire                                        std__mgr14__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane7_strm0_data        ,
            output  wire                                        mgr14__std__lane7_strm0_data_valid  ,

            // manager 14, lane 7, stream 1      
            input   wire                                        std__mgr14__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane7_strm1_data        ,
            output  wire                                        mgr14__std__lane7_strm1_data_valid  ,

            // manager 14, lane 8, stream 0      
            input   wire                                        std__mgr14__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane8_strm0_data        ,
            output  wire                                        mgr14__std__lane8_strm0_data_valid  ,

            // manager 14, lane 8, stream 1      
            input   wire                                        std__mgr14__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane8_strm1_data        ,
            output  wire                                        mgr14__std__lane8_strm1_data_valid  ,

            // manager 14, lane 9, stream 0      
            input   wire                                        std__mgr14__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane9_strm0_data        ,
            output  wire                                        mgr14__std__lane9_strm0_data_valid  ,

            // manager 14, lane 9, stream 1      
            input   wire                                        std__mgr14__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane9_strm1_data        ,
            output  wire                                        mgr14__std__lane9_strm1_data_valid  ,

            // manager 14, lane 10, stream 0      
            input   wire                                        std__mgr14__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane10_strm0_data        ,
            output  wire                                        mgr14__std__lane10_strm0_data_valid  ,

            // manager 14, lane 10, stream 1      
            input   wire                                        std__mgr14__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane10_strm1_data        ,
            output  wire                                        mgr14__std__lane10_strm1_data_valid  ,

            // manager 14, lane 11, stream 0      
            input   wire                                        std__mgr14__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane11_strm0_data        ,
            output  wire                                        mgr14__std__lane11_strm0_data_valid  ,

            // manager 14, lane 11, stream 1      
            input   wire                                        std__mgr14__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane11_strm1_data        ,
            output  wire                                        mgr14__std__lane11_strm1_data_valid  ,

            // manager 14, lane 12, stream 0      
            input   wire                                        std__mgr14__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane12_strm0_data        ,
            output  wire                                        mgr14__std__lane12_strm0_data_valid  ,

            // manager 14, lane 12, stream 1      
            input   wire                                        std__mgr14__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane12_strm1_data        ,
            output  wire                                        mgr14__std__lane12_strm1_data_valid  ,

            // manager 14, lane 13, stream 0      
            input   wire                                        std__mgr14__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane13_strm0_data        ,
            output  wire                                        mgr14__std__lane13_strm0_data_valid  ,

            // manager 14, lane 13, stream 1      
            input   wire                                        std__mgr14__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane13_strm1_data        ,
            output  wire                                        mgr14__std__lane13_strm1_data_valid  ,

            // manager 14, lane 14, stream 0      
            input   wire                                        std__mgr14__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane14_strm0_data        ,
            output  wire                                        mgr14__std__lane14_strm0_data_valid  ,

            // manager 14, lane 14, stream 1      
            input   wire                                        std__mgr14__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane14_strm1_data        ,
            output  wire                                        mgr14__std__lane14_strm1_data_valid  ,

            // manager 14, lane 15, stream 0      
            input   wire                                        std__mgr14__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane15_strm0_data        ,
            output  wire                                        mgr14__std__lane15_strm0_data_valid  ,

            // manager 14, lane 15, stream 1      
            input   wire                                        std__mgr14__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane15_strm1_data        ,
            output  wire                                        mgr14__std__lane15_strm1_data_valid  ,

            // manager 14, lane 16, stream 0      
            input   wire                                        std__mgr14__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane16_strm0_data        ,
            output  wire                                        mgr14__std__lane16_strm0_data_valid  ,

            // manager 14, lane 16, stream 1      
            input   wire                                        std__mgr14__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane16_strm1_data        ,
            output  wire                                        mgr14__std__lane16_strm1_data_valid  ,

            // manager 14, lane 17, stream 0      
            input   wire                                        std__mgr14__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane17_strm0_data        ,
            output  wire                                        mgr14__std__lane17_strm0_data_valid  ,

            // manager 14, lane 17, stream 1      
            input   wire                                        std__mgr14__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane17_strm1_data        ,
            output  wire                                        mgr14__std__lane17_strm1_data_valid  ,

            // manager 14, lane 18, stream 0      
            input   wire                                        std__mgr14__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane18_strm0_data        ,
            output  wire                                        mgr14__std__lane18_strm0_data_valid  ,

            // manager 14, lane 18, stream 1      
            input   wire                                        std__mgr14__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane18_strm1_data        ,
            output  wire                                        mgr14__std__lane18_strm1_data_valid  ,

            // manager 14, lane 19, stream 0      
            input   wire                                        std__mgr14__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane19_strm0_data        ,
            output  wire                                        mgr14__std__lane19_strm0_data_valid  ,

            // manager 14, lane 19, stream 1      
            input   wire                                        std__mgr14__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane19_strm1_data        ,
            output  wire                                        mgr14__std__lane19_strm1_data_valid  ,

            // manager 14, lane 20, stream 0      
            input   wire                                        std__mgr14__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane20_strm0_data        ,
            output  wire                                        mgr14__std__lane20_strm0_data_valid  ,

            // manager 14, lane 20, stream 1      
            input   wire                                        std__mgr14__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane20_strm1_data        ,
            output  wire                                        mgr14__std__lane20_strm1_data_valid  ,

            // manager 14, lane 21, stream 0      
            input   wire                                        std__mgr14__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane21_strm0_data        ,
            output  wire                                        mgr14__std__lane21_strm0_data_valid  ,

            // manager 14, lane 21, stream 1      
            input   wire                                        std__mgr14__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane21_strm1_data        ,
            output  wire                                        mgr14__std__lane21_strm1_data_valid  ,

            // manager 14, lane 22, stream 0      
            input   wire                                        std__mgr14__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane22_strm0_data        ,
            output  wire                                        mgr14__std__lane22_strm0_data_valid  ,

            // manager 14, lane 22, stream 1      
            input   wire                                        std__mgr14__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane22_strm1_data        ,
            output  wire                                        mgr14__std__lane22_strm1_data_valid  ,

            // manager 14, lane 23, stream 0      
            input   wire                                        std__mgr14__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane23_strm0_data        ,
            output  wire                                        mgr14__std__lane23_strm0_data_valid  ,

            // manager 14, lane 23, stream 1      
            input   wire                                        std__mgr14__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane23_strm1_data        ,
            output  wire                                        mgr14__std__lane23_strm1_data_valid  ,

            // manager 14, lane 24, stream 0      
            input   wire                                        std__mgr14__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane24_strm0_data        ,
            output  wire                                        mgr14__std__lane24_strm0_data_valid  ,

            // manager 14, lane 24, stream 1      
            input   wire                                        std__mgr14__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane24_strm1_data        ,
            output  wire                                        mgr14__std__lane24_strm1_data_valid  ,

            // manager 14, lane 25, stream 0      
            input   wire                                        std__mgr14__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane25_strm0_data        ,
            output  wire                                        mgr14__std__lane25_strm0_data_valid  ,

            // manager 14, lane 25, stream 1      
            input   wire                                        std__mgr14__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane25_strm1_data        ,
            output  wire                                        mgr14__std__lane25_strm1_data_valid  ,

            // manager 14, lane 26, stream 0      
            input   wire                                        std__mgr14__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane26_strm0_data        ,
            output  wire                                        mgr14__std__lane26_strm0_data_valid  ,

            // manager 14, lane 26, stream 1      
            input   wire                                        std__mgr14__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane26_strm1_data        ,
            output  wire                                        mgr14__std__lane26_strm1_data_valid  ,

            // manager 14, lane 27, stream 0      
            input   wire                                        std__mgr14__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane27_strm0_data        ,
            output  wire                                        mgr14__std__lane27_strm0_data_valid  ,

            // manager 14, lane 27, stream 1      
            input   wire                                        std__mgr14__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane27_strm1_data        ,
            output  wire                                        mgr14__std__lane27_strm1_data_valid  ,

            // manager 14, lane 28, stream 0      
            input   wire                                        std__mgr14__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane28_strm0_data        ,
            output  wire                                        mgr14__std__lane28_strm0_data_valid  ,

            // manager 14, lane 28, stream 1      
            input   wire                                        std__mgr14__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane28_strm1_data        ,
            output  wire                                        mgr14__std__lane28_strm1_data_valid  ,

            // manager 14, lane 29, stream 0      
            input   wire                                        std__mgr14__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane29_strm0_data        ,
            output  wire                                        mgr14__std__lane29_strm0_data_valid  ,

            // manager 14, lane 29, stream 1      
            input   wire                                        std__mgr14__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane29_strm1_data        ,
            output  wire                                        mgr14__std__lane29_strm1_data_valid  ,

            // manager 14, lane 30, stream 0      
            input   wire                                        std__mgr14__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane30_strm0_data        ,
            output  wire                                        mgr14__std__lane30_strm0_data_valid  ,

            // manager 14, lane 30, stream 1      
            input   wire                                        std__mgr14__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane30_strm1_data        ,
            output  wire                                        mgr14__std__lane30_strm1_data_valid  ,

            // manager 14, lane 31, stream 0      
            input   wire                                        std__mgr14__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane31_strm0_data        ,
            output  wire                                        mgr14__std__lane31_strm0_data_valid  ,

            // manager 14, lane 31, stream 1      
            input   wire                                        std__mgr14__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr14__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr14__std__lane31_strm1_data        ,
            output  wire                                        mgr14__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 15, lane 0, stream 0      
            input   wire                                        std__mgr15__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane0_strm0_data        ,
            output  wire                                        mgr15__std__lane0_strm0_data_valid  ,

            // manager 15, lane 0, stream 1      
            input   wire                                        std__mgr15__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane0_strm1_data        ,
            output  wire                                        mgr15__std__lane0_strm1_data_valid  ,

            // manager 15, lane 1, stream 0      
            input   wire                                        std__mgr15__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane1_strm0_data        ,
            output  wire                                        mgr15__std__lane1_strm0_data_valid  ,

            // manager 15, lane 1, stream 1      
            input   wire                                        std__mgr15__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane1_strm1_data        ,
            output  wire                                        mgr15__std__lane1_strm1_data_valid  ,

            // manager 15, lane 2, stream 0      
            input   wire                                        std__mgr15__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane2_strm0_data        ,
            output  wire                                        mgr15__std__lane2_strm0_data_valid  ,

            // manager 15, lane 2, stream 1      
            input   wire                                        std__mgr15__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane2_strm1_data        ,
            output  wire                                        mgr15__std__lane2_strm1_data_valid  ,

            // manager 15, lane 3, stream 0      
            input   wire                                        std__mgr15__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane3_strm0_data        ,
            output  wire                                        mgr15__std__lane3_strm0_data_valid  ,

            // manager 15, lane 3, stream 1      
            input   wire                                        std__mgr15__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane3_strm1_data        ,
            output  wire                                        mgr15__std__lane3_strm1_data_valid  ,

            // manager 15, lane 4, stream 0      
            input   wire                                        std__mgr15__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane4_strm0_data        ,
            output  wire                                        mgr15__std__lane4_strm0_data_valid  ,

            // manager 15, lane 4, stream 1      
            input   wire                                        std__mgr15__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane4_strm1_data        ,
            output  wire                                        mgr15__std__lane4_strm1_data_valid  ,

            // manager 15, lane 5, stream 0      
            input   wire                                        std__mgr15__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane5_strm0_data        ,
            output  wire                                        mgr15__std__lane5_strm0_data_valid  ,

            // manager 15, lane 5, stream 1      
            input   wire                                        std__mgr15__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane5_strm1_data        ,
            output  wire                                        mgr15__std__lane5_strm1_data_valid  ,

            // manager 15, lane 6, stream 0      
            input   wire                                        std__mgr15__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane6_strm0_data        ,
            output  wire                                        mgr15__std__lane6_strm0_data_valid  ,

            // manager 15, lane 6, stream 1      
            input   wire                                        std__mgr15__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane6_strm1_data        ,
            output  wire                                        mgr15__std__lane6_strm1_data_valid  ,

            // manager 15, lane 7, stream 0      
            input   wire                                        std__mgr15__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane7_strm0_data        ,
            output  wire                                        mgr15__std__lane7_strm0_data_valid  ,

            // manager 15, lane 7, stream 1      
            input   wire                                        std__mgr15__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane7_strm1_data        ,
            output  wire                                        mgr15__std__lane7_strm1_data_valid  ,

            // manager 15, lane 8, stream 0      
            input   wire                                        std__mgr15__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane8_strm0_data        ,
            output  wire                                        mgr15__std__lane8_strm0_data_valid  ,

            // manager 15, lane 8, stream 1      
            input   wire                                        std__mgr15__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane8_strm1_data        ,
            output  wire                                        mgr15__std__lane8_strm1_data_valid  ,

            // manager 15, lane 9, stream 0      
            input   wire                                        std__mgr15__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane9_strm0_data        ,
            output  wire                                        mgr15__std__lane9_strm0_data_valid  ,

            // manager 15, lane 9, stream 1      
            input   wire                                        std__mgr15__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane9_strm1_data        ,
            output  wire                                        mgr15__std__lane9_strm1_data_valid  ,

            // manager 15, lane 10, stream 0      
            input   wire                                        std__mgr15__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane10_strm0_data        ,
            output  wire                                        mgr15__std__lane10_strm0_data_valid  ,

            // manager 15, lane 10, stream 1      
            input   wire                                        std__mgr15__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane10_strm1_data        ,
            output  wire                                        mgr15__std__lane10_strm1_data_valid  ,

            // manager 15, lane 11, stream 0      
            input   wire                                        std__mgr15__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane11_strm0_data        ,
            output  wire                                        mgr15__std__lane11_strm0_data_valid  ,

            // manager 15, lane 11, stream 1      
            input   wire                                        std__mgr15__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane11_strm1_data        ,
            output  wire                                        mgr15__std__lane11_strm1_data_valid  ,

            // manager 15, lane 12, stream 0      
            input   wire                                        std__mgr15__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane12_strm0_data        ,
            output  wire                                        mgr15__std__lane12_strm0_data_valid  ,

            // manager 15, lane 12, stream 1      
            input   wire                                        std__mgr15__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane12_strm1_data        ,
            output  wire                                        mgr15__std__lane12_strm1_data_valid  ,

            // manager 15, lane 13, stream 0      
            input   wire                                        std__mgr15__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane13_strm0_data        ,
            output  wire                                        mgr15__std__lane13_strm0_data_valid  ,

            // manager 15, lane 13, stream 1      
            input   wire                                        std__mgr15__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane13_strm1_data        ,
            output  wire                                        mgr15__std__lane13_strm1_data_valid  ,

            // manager 15, lane 14, stream 0      
            input   wire                                        std__mgr15__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane14_strm0_data        ,
            output  wire                                        mgr15__std__lane14_strm0_data_valid  ,

            // manager 15, lane 14, stream 1      
            input   wire                                        std__mgr15__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane14_strm1_data        ,
            output  wire                                        mgr15__std__lane14_strm1_data_valid  ,

            // manager 15, lane 15, stream 0      
            input   wire                                        std__mgr15__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane15_strm0_data        ,
            output  wire                                        mgr15__std__lane15_strm0_data_valid  ,

            // manager 15, lane 15, stream 1      
            input   wire                                        std__mgr15__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane15_strm1_data        ,
            output  wire                                        mgr15__std__lane15_strm1_data_valid  ,

            // manager 15, lane 16, stream 0      
            input   wire                                        std__mgr15__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane16_strm0_data        ,
            output  wire                                        mgr15__std__lane16_strm0_data_valid  ,

            // manager 15, lane 16, stream 1      
            input   wire                                        std__mgr15__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane16_strm1_data        ,
            output  wire                                        mgr15__std__lane16_strm1_data_valid  ,

            // manager 15, lane 17, stream 0      
            input   wire                                        std__mgr15__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane17_strm0_data        ,
            output  wire                                        mgr15__std__lane17_strm0_data_valid  ,

            // manager 15, lane 17, stream 1      
            input   wire                                        std__mgr15__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane17_strm1_data        ,
            output  wire                                        mgr15__std__lane17_strm1_data_valid  ,

            // manager 15, lane 18, stream 0      
            input   wire                                        std__mgr15__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane18_strm0_data        ,
            output  wire                                        mgr15__std__lane18_strm0_data_valid  ,

            // manager 15, lane 18, stream 1      
            input   wire                                        std__mgr15__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane18_strm1_data        ,
            output  wire                                        mgr15__std__lane18_strm1_data_valid  ,

            // manager 15, lane 19, stream 0      
            input   wire                                        std__mgr15__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane19_strm0_data        ,
            output  wire                                        mgr15__std__lane19_strm0_data_valid  ,

            // manager 15, lane 19, stream 1      
            input   wire                                        std__mgr15__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane19_strm1_data        ,
            output  wire                                        mgr15__std__lane19_strm1_data_valid  ,

            // manager 15, lane 20, stream 0      
            input   wire                                        std__mgr15__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane20_strm0_data        ,
            output  wire                                        mgr15__std__lane20_strm0_data_valid  ,

            // manager 15, lane 20, stream 1      
            input   wire                                        std__mgr15__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane20_strm1_data        ,
            output  wire                                        mgr15__std__lane20_strm1_data_valid  ,

            // manager 15, lane 21, stream 0      
            input   wire                                        std__mgr15__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane21_strm0_data        ,
            output  wire                                        mgr15__std__lane21_strm0_data_valid  ,

            // manager 15, lane 21, stream 1      
            input   wire                                        std__mgr15__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane21_strm1_data        ,
            output  wire                                        mgr15__std__lane21_strm1_data_valid  ,

            // manager 15, lane 22, stream 0      
            input   wire                                        std__mgr15__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane22_strm0_data        ,
            output  wire                                        mgr15__std__lane22_strm0_data_valid  ,

            // manager 15, lane 22, stream 1      
            input   wire                                        std__mgr15__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane22_strm1_data        ,
            output  wire                                        mgr15__std__lane22_strm1_data_valid  ,

            // manager 15, lane 23, stream 0      
            input   wire                                        std__mgr15__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane23_strm0_data        ,
            output  wire                                        mgr15__std__lane23_strm0_data_valid  ,

            // manager 15, lane 23, stream 1      
            input   wire                                        std__mgr15__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane23_strm1_data        ,
            output  wire                                        mgr15__std__lane23_strm1_data_valid  ,

            // manager 15, lane 24, stream 0      
            input   wire                                        std__mgr15__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane24_strm0_data        ,
            output  wire                                        mgr15__std__lane24_strm0_data_valid  ,

            // manager 15, lane 24, stream 1      
            input   wire                                        std__mgr15__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane24_strm1_data        ,
            output  wire                                        mgr15__std__lane24_strm1_data_valid  ,

            // manager 15, lane 25, stream 0      
            input   wire                                        std__mgr15__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane25_strm0_data        ,
            output  wire                                        mgr15__std__lane25_strm0_data_valid  ,

            // manager 15, lane 25, stream 1      
            input   wire                                        std__mgr15__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane25_strm1_data        ,
            output  wire                                        mgr15__std__lane25_strm1_data_valid  ,

            // manager 15, lane 26, stream 0      
            input   wire                                        std__mgr15__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane26_strm0_data        ,
            output  wire                                        mgr15__std__lane26_strm0_data_valid  ,

            // manager 15, lane 26, stream 1      
            input   wire                                        std__mgr15__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane26_strm1_data        ,
            output  wire                                        mgr15__std__lane26_strm1_data_valid  ,

            // manager 15, lane 27, stream 0      
            input   wire                                        std__mgr15__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane27_strm0_data        ,
            output  wire                                        mgr15__std__lane27_strm0_data_valid  ,

            // manager 15, lane 27, stream 1      
            input   wire                                        std__mgr15__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane27_strm1_data        ,
            output  wire                                        mgr15__std__lane27_strm1_data_valid  ,

            // manager 15, lane 28, stream 0      
            input   wire                                        std__mgr15__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane28_strm0_data        ,
            output  wire                                        mgr15__std__lane28_strm0_data_valid  ,

            // manager 15, lane 28, stream 1      
            input   wire                                        std__mgr15__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane28_strm1_data        ,
            output  wire                                        mgr15__std__lane28_strm1_data_valid  ,

            // manager 15, lane 29, stream 0      
            input   wire                                        std__mgr15__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane29_strm0_data        ,
            output  wire                                        mgr15__std__lane29_strm0_data_valid  ,

            // manager 15, lane 29, stream 1      
            input   wire                                        std__mgr15__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane29_strm1_data        ,
            output  wire                                        mgr15__std__lane29_strm1_data_valid  ,

            // manager 15, lane 30, stream 0      
            input   wire                                        std__mgr15__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane30_strm0_data        ,
            output  wire                                        mgr15__std__lane30_strm0_data_valid  ,

            // manager 15, lane 30, stream 1      
            input   wire                                        std__mgr15__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane30_strm1_data        ,
            output  wire                                        mgr15__std__lane30_strm1_data_valid  ,

            // manager 15, lane 31, stream 0      
            input   wire                                        std__mgr15__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane31_strm0_data        ,
            output  wire                                        mgr15__std__lane31_strm0_data_valid  ,

            // manager 15, lane 31, stream 1      
            input   wire                                        std__mgr15__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr15__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr15__std__lane31_strm1_data        ,
            output  wire                                        mgr15__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 16, lane 0, stream 0      
            input   wire                                        std__mgr16__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane0_strm0_data        ,
            output  wire                                        mgr16__std__lane0_strm0_data_valid  ,

            // manager 16, lane 0, stream 1      
            input   wire                                        std__mgr16__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane0_strm1_data        ,
            output  wire                                        mgr16__std__lane0_strm1_data_valid  ,

            // manager 16, lane 1, stream 0      
            input   wire                                        std__mgr16__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane1_strm0_data        ,
            output  wire                                        mgr16__std__lane1_strm0_data_valid  ,

            // manager 16, lane 1, stream 1      
            input   wire                                        std__mgr16__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane1_strm1_data        ,
            output  wire                                        mgr16__std__lane1_strm1_data_valid  ,

            // manager 16, lane 2, stream 0      
            input   wire                                        std__mgr16__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane2_strm0_data        ,
            output  wire                                        mgr16__std__lane2_strm0_data_valid  ,

            // manager 16, lane 2, stream 1      
            input   wire                                        std__mgr16__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane2_strm1_data        ,
            output  wire                                        mgr16__std__lane2_strm1_data_valid  ,

            // manager 16, lane 3, stream 0      
            input   wire                                        std__mgr16__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane3_strm0_data        ,
            output  wire                                        mgr16__std__lane3_strm0_data_valid  ,

            // manager 16, lane 3, stream 1      
            input   wire                                        std__mgr16__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane3_strm1_data        ,
            output  wire                                        mgr16__std__lane3_strm1_data_valid  ,

            // manager 16, lane 4, stream 0      
            input   wire                                        std__mgr16__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane4_strm0_data        ,
            output  wire                                        mgr16__std__lane4_strm0_data_valid  ,

            // manager 16, lane 4, stream 1      
            input   wire                                        std__mgr16__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane4_strm1_data        ,
            output  wire                                        mgr16__std__lane4_strm1_data_valid  ,

            // manager 16, lane 5, stream 0      
            input   wire                                        std__mgr16__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane5_strm0_data        ,
            output  wire                                        mgr16__std__lane5_strm0_data_valid  ,

            // manager 16, lane 5, stream 1      
            input   wire                                        std__mgr16__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane5_strm1_data        ,
            output  wire                                        mgr16__std__lane5_strm1_data_valid  ,

            // manager 16, lane 6, stream 0      
            input   wire                                        std__mgr16__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane6_strm0_data        ,
            output  wire                                        mgr16__std__lane6_strm0_data_valid  ,

            // manager 16, lane 6, stream 1      
            input   wire                                        std__mgr16__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane6_strm1_data        ,
            output  wire                                        mgr16__std__lane6_strm1_data_valid  ,

            // manager 16, lane 7, stream 0      
            input   wire                                        std__mgr16__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane7_strm0_data        ,
            output  wire                                        mgr16__std__lane7_strm0_data_valid  ,

            // manager 16, lane 7, stream 1      
            input   wire                                        std__mgr16__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane7_strm1_data        ,
            output  wire                                        mgr16__std__lane7_strm1_data_valid  ,

            // manager 16, lane 8, stream 0      
            input   wire                                        std__mgr16__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane8_strm0_data        ,
            output  wire                                        mgr16__std__lane8_strm0_data_valid  ,

            // manager 16, lane 8, stream 1      
            input   wire                                        std__mgr16__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane8_strm1_data        ,
            output  wire                                        mgr16__std__lane8_strm1_data_valid  ,

            // manager 16, lane 9, stream 0      
            input   wire                                        std__mgr16__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane9_strm0_data        ,
            output  wire                                        mgr16__std__lane9_strm0_data_valid  ,

            // manager 16, lane 9, stream 1      
            input   wire                                        std__mgr16__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane9_strm1_data        ,
            output  wire                                        mgr16__std__lane9_strm1_data_valid  ,

            // manager 16, lane 10, stream 0      
            input   wire                                        std__mgr16__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane10_strm0_data        ,
            output  wire                                        mgr16__std__lane10_strm0_data_valid  ,

            // manager 16, lane 10, stream 1      
            input   wire                                        std__mgr16__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane10_strm1_data        ,
            output  wire                                        mgr16__std__lane10_strm1_data_valid  ,

            // manager 16, lane 11, stream 0      
            input   wire                                        std__mgr16__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane11_strm0_data        ,
            output  wire                                        mgr16__std__lane11_strm0_data_valid  ,

            // manager 16, lane 11, stream 1      
            input   wire                                        std__mgr16__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane11_strm1_data        ,
            output  wire                                        mgr16__std__lane11_strm1_data_valid  ,

            // manager 16, lane 12, stream 0      
            input   wire                                        std__mgr16__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane12_strm0_data        ,
            output  wire                                        mgr16__std__lane12_strm0_data_valid  ,

            // manager 16, lane 12, stream 1      
            input   wire                                        std__mgr16__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane12_strm1_data        ,
            output  wire                                        mgr16__std__lane12_strm1_data_valid  ,

            // manager 16, lane 13, stream 0      
            input   wire                                        std__mgr16__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane13_strm0_data        ,
            output  wire                                        mgr16__std__lane13_strm0_data_valid  ,

            // manager 16, lane 13, stream 1      
            input   wire                                        std__mgr16__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane13_strm1_data        ,
            output  wire                                        mgr16__std__lane13_strm1_data_valid  ,

            // manager 16, lane 14, stream 0      
            input   wire                                        std__mgr16__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane14_strm0_data        ,
            output  wire                                        mgr16__std__lane14_strm0_data_valid  ,

            // manager 16, lane 14, stream 1      
            input   wire                                        std__mgr16__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane14_strm1_data        ,
            output  wire                                        mgr16__std__lane14_strm1_data_valid  ,

            // manager 16, lane 15, stream 0      
            input   wire                                        std__mgr16__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane15_strm0_data        ,
            output  wire                                        mgr16__std__lane15_strm0_data_valid  ,

            // manager 16, lane 15, stream 1      
            input   wire                                        std__mgr16__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane15_strm1_data        ,
            output  wire                                        mgr16__std__lane15_strm1_data_valid  ,

            // manager 16, lane 16, stream 0      
            input   wire                                        std__mgr16__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane16_strm0_data        ,
            output  wire                                        mgr16__std__lane16_strm0_data_valid  ,

            // manager 16, lane 16, stream 1      
            input   wire                                        std__mgr16__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane16_strm1_data        ,
            output  wire                                        mgr16__std__lane16_strm1_data_valid  ,

            // manager 16, lane 17, stream 0      
            input   wire                                        std__mgr16__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane17_strm0_data        ,
            output  wire                                        mgr16__std__lane17_strm0_data_valid  ,

            // manager 16, lane 17, stream 1      
            input   wire                                        std__mgr16__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane17_strm1_data        ,
            output  wire                                        mgr16__std__lane17_strm1_data_valid  ,

            // manager 16, lane 18, stream 0      
            input   wire                                        std__mgr16__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane18_strm0_data        ,
            output  wire                                        mgr16__std__lane18_strm0_data_valid  ,

            // manager 16, lane 18, stream 1      
            input   wire                                        std__mgr16__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane18_strm1_data        ,
            output  wire                                        mgr16__std__lane18_strm1_data_valid  ,

            // manager 16, lane 19, stream 0      
            input   wire                                        std__mgr16__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane19_strm0_data        ,
            output  wire                                        mgr16__std__lane19_strm0_data_valid  ,

            // manager 16, lane 19, stream 1      
            input   wire                                        std__mgr16__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane19_strm1_data        ,
            output  wire                                        mgr16__std__lane19_strm1_data_valid  ,

            // manager 16, lane 20, stream 0      
            input   wire                                        std__mgr16__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane20_strm0_data        ,
            output  wire                                        mgr16__std__lane20_strm0_data_valid  ,

            // manager 16, lane 20, stream 1      
            input   wire                                        std__mgr16__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane20_strm1_data        ,
            output  wire                                        mgr16__std__lane20_strm1_data_valid  ,

            // manager 16, lane 21, stream 0      
            input   wire                                        std__mgr16__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane21_strm0_data        ,
            output  wire                                        mgr16__std__lane21_strm0_data_valid  ,

            // manager 16, lane 21, stream 1      
            input   wire                                        std__mgr16__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane21_strm1_data        ,
            output  wire                                        mgr16__std__lane21_strm1_data_valid  ,

            // manager 16, lane 22, stream 0      
            input   wire                                        std__mgr16__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane22_strm0_data        ,
            output  wire                                        mgr16__std__lane22_strm0_data_valid  ,

            // manager 16, lane 22, stream 1      
            input   wire                                        std__mgr16__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane22_strm1_data        ,
            output  wire                                        mgr16__std__lane22_strm1_data_valid  ,

            // manager 16, lane 23, stream 0      
            input   wire                                        std__mgr16__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane23_strm0_data        ,
            output  wire                                        mgr16__std__lane23_strm0_data_valid  ,

            // manager 16, lane 23, stream 1      
            input   wire                                        std__mgr16__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane23_strm1_data        ,
            output  wire                                        mgr16__std__lane23_strm1_data_valid  ,

            // manager 16, lane 24, stream 0      
            input   wire                                        std__mgr16__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane24_strm0_data        ,
            output  wire                                        mgr16__std__lane24_strm0_data_valid  ,

            // manager 16, lane 24, stream 1      
            input   wire                                        std__mgr16__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane24_strm1_data        ,
            output  wire                                        mgr16__std__lane24_strm1_data_valid  ,

            // manager 16, lane 25, stream 0      
            input   wire                                        std__mgr16__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane25_strm0_data        ,
            output  wire                                        mgr16__std__lane25_strm0_data_valid  ,

            // manager 16, lane 25, stream 1      
            input   wire                                        std__mgr16__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane25_strm1_data        ,
            output  wire                                        mgr16__std__lane25_strm1_data_valid  ,

            // manager 16, lane 26, stream 0      
            input   wire                                        std__mgr16__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane26_strm0_data        ,
            output  wire                                        mgr16__std__lane26_strm0_data_valid  ,

            // manager 16, lane 26, stream 1      
            input   wire                                        std__mgr16__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane26_strm1_data        ,
            output  wire                                        mgr16__std__lane26_strm1_data_valid  ,

            // manager 16, lane 27, stream 0      
            input   wire                                        std__mgr16__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane27_strm0_data        ,
            output  wire                                        mgr16__std__lane27_strm0_data_valid  ,

            // manager 16, lane 27, stream 1      
            input   wire                                        std__mgr16__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane27_strm1_data        ,
            output  wire                                        mgr16__std__lane27_strm1_data_valid  ,

            // manager 16, lane 28, stream 0      
            input   wire                                        std__mgr16__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane28_strm0_data        ,
            output  wire                                        mgr16__std__lane28_strm0_data_valid  ,

            // manager 16, lane 28, stream 1      
            input   wire                                        std__mgr16__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane28_strm1_data        ,
            output  wire                                        mgr16__std__lane28_strm1_data_valid  ,

            // manager 16, lane 29, stream 0      
            input   wire                                        std__mgr16__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane29_strm0_data        ,
            output  wire                                        mgr16__std__lane29_strm0_data_valid  ,

            // manager 16, lane 29, stream 1      
            input   wire                                        std__mgr16__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane29_strm1_data        ,
            output  wire                                        mgr16__std__lane29_strm1_data_valid  ,

            // manager 16, lane 30, stream 0      
            input   wire                                        std__mgr16__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane30_strm0_data        ,
            output  wire                                        mgr16__std__lane30_strm0_data_valid  ,

            // manager 16, lane 30, stream 1      
            input   wire                                        std__mgr16__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane30_strm1_data        ,
            output  wire                                        mgr16__std__lane30_strm1_data_valid  ,

            // manager 16, lane 31, stream 0      
            input   wire                                        std__mgr16__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane31_strm0_data        ,
            output  wire                                        mgr16__std__lane31_strm0_data_valid  ,

            // manager 16, lane 31, stream 1      
            input   wire                                        std__mgr16__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr16__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr16__std__lane31_strm1_data        ,
            output  wire                                        mgr16__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 17, lane 0, stream 0      
            input   wire                                        std__mgr17__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane0_strm0_data        ,
            output  wire                                        mgr17__std__lane0_strm0_data_valid  ,

            // manager 17, lane 0, stream 1      
            input   wire                                        std__mgr17__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane0_strm1_data        ,
            output  wire                                        mgr17__std__lane0_strm1_data_valid  ,

            // manager 17, lane 1, stream 0      
            input   wire                                        std__mgr17__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane1_strm0_data        ,
            output  wire                                        mgr17__std__lane1_strm0_data_valid  ,

            // manager 17, lane 1, stream 1      
            input   wire                                        std__mgr17__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane1_strm1_data        ,
            output  wire                                        mgr17__std__lane1_strm1_data_valid  ,

            // manager 17, lane 2, stream 0      
            input   wire                                        std__mgr17__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane2_strm0_data        ,
            output  wire                                        mgr17__std__lane2_strm0_data_valid  ,

            // manager 17, lane 2, stream 1      
            input   wire                                        std__mgr17__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane2_strm1_data        ,
            output  wire                                        mgr17__std__lane2_strm1_data_valid  ,

            // manager 17, lane 3, stream 0      
            input   wire                                        std__mgr17__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane3_strm0_data        ,
            output  wire                                        mgr17__std__lane3_strm0_data_valid  ,

            // manager 17, lane 3, stream 1      
            input   wire                                        std__mgr17__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane3_strm1_data        ,
            output  wire                                        mgr17__std__lane3_strm1_data_valid  ,

            // manager 17, lane 4, stream 0      
            input   wire                                        std__mgr17__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane4_strm0_data        ,
            output  wire                                        mgr17__std__lane4_strm0_data_valid  ,

            // manager 17, lane 4, stream 1      
            input   wire                                        std__mgr17__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane4_strm1_data        ,
            output  wire                                        mgr17__std__lane4_strm1_data_valid  ,

            // manager 17, lane 5, stream 0      
            input   wire                                        std__mgr17__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane5_strm0_data        ,
            output  wire                                        mgr17__std__lane5_strm0_data_valid  ,

            // manager 17, lane 5, stream 1      
            input   wire                                        std__mgr17__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane5_strm1_data        ,
            output  wire                                        mgr17__std__lane5_strm1_data_valid  ,

            // manager 17, lane 6, stream 0      
            input   wire                                        std__mgr17__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane6_strm0_data        ,
            output  wire                                        mgr17__std__lane6_strm0_data_valid  ,

            // manager 17, lane 6, stream 1      
            input   wire                                        std__mgr17__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane6_strm1_data        ,
            output  wire                                        mgr17__std__lane6_strm1_data_valid  ,

            // manager 17, lane 7, stream 0      
            input   wire                                        std__mgr17__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane7_strm0_data        ,
            output  wire                                        mgr17__std__lane7_strm0_data_valid  ,

            // manager 17, lane 7, stream 1      
            input   wire                                        std__mgr17__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane7_strm1_data        ,
            output  wire                                        mgr17__std__lane7_strm1_data_valid  ,

            // manager 17, lane 8, stream 0      
            input   wire                                        std__mgr17__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane8_strm0_data        ,
            output  wire                                        mgr17__std__lane8_strm0_data_valid  ,

            // manager 17, lane 8, stream 1      
            input   wire                                        std__mgr17__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane8_strm1_data        ,
            output  wire                                        mgr17__std__lane8_strm1_data_valid  ,

            // manager 17, lane 9, stream 0      
            input   wire                                        std__mgr17__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane9_strm0_data        ,
            output  wire                                        mgr17__std__lane9_strm0_data_valid  ,

            // manager 17, lane 9, stream 1      
            input   wire                                        std__mgr17__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane9_strm1_data        ,
            output  wire                                        mgr17__std__lane9_strm1_data_valid  ,

            // manager 17, lane 10, stream 0      
            input   wire                                        std__mgr17__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane10_strm0_data        ,
            output  wire                                        mgr17__std__lane10_strm0_data_valid  ,

            // manager 17, lane 10, stream 1      
            input   wire                                        std__mgr17__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane10_strm1_data        ,
            output  wire                                        mgr17__std__lane10_strm1_data_valid  ,

            // manager 17, lane 11, stream 0      
            input   wire                                        std__mgr17__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane11_strm0_data        ,
            output  wire                                        mgr17__std__lane11_strm0_data_valid  ,

            // manager 17, lane 11, stream 1      
            input   wire                                        std__mgr17__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane11_strm1_data        ,
            output  wire                                        mgr17__std__lane11_strm1_data_valid  ,

            // manager 17, lane 12, stream 0      
            input   wire                                        std__mgr17__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane12_strm0_data        ,
            output  wire                                        mgr17__std__lane12_strm0_data_valid  ,

            // manager 17, lane 12, stream 1      
            input   wire                                        std__mgr17__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane12_strm1_data        ,
            output  wire                                        mgr17__std__lane12_strm1_data_valid  ,

            // manager 17, lane 13, stream 0      
            input   wire                                        std__mgr17__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane13_strm0_data        ,
            output  wire                                        mgr17__std__lane13_strm0_data_valid  ,

            // manager 17, lane 13, stream 1      
            input   wire                                        std__mgr17__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane13_strm1_data        ,
            output  wire                                        mgr17__std__lane13_strm1_data_valid  ,

            // manager 17, lane 14, stream 0      
            input   wire                                        std__mgr17__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane14_strm0_data        ,
            output  wire                                        mgr17__std__lane14_strm0_data_valid  ,

            // manager 17, lane 14, stream 1      
            input   wire                                        std__mgr17__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane14_strm1_data        ,
            output  wire                                        mgr17__std__lane14_strm1_data_valid  ,

            // manager 17, lane 15, stream 0      
            input   wire                                        std__mgr17__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane15_strm0_data        ,
            output  wire                                        mgr17__std__lane15_strm0_data_valid  ,

            // manager 17, lane 15, stream 1      
            input   wire                                        std__mgr17__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane15_strm1_data        ,
            output  wire                                        mgr17__std__lane15_strm1_data_valid  ,

            // manager 17, lane 16, stream 0      
            input   wire                                        std__mgr17__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane16_strm0_data        ,
            output  wire                                        mgr17__std__lane16_strm0_data_valid  ,

            // manager 17, lane 16, stream 1      
            input   wire                                        std__mgr17__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane16_strm1_data        ,
            output  wire                                        mgr17__std__lane16_strm1_data_valid  ,

            // manager 17, lane 17, stream 0      
            input   wire                                        std__mgr17__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane17_strm0_data        ,
            output  wire                                        mgr17__std__lane17_strm0_data_valid  ,

            // manager 17, lane 17, stream 1      
            input   wire                                        std__mgr17__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane17_strm1_data        ,
            output  wire                                        mgr17__std__lane17_strm1_data_valid  ,

            // manager 17, lane 18, stream 0      
            input   wire                                        std__mgr17__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane18_strm0_data        ,
            output  wire                                        mgr17__std__lane18_strm0_data_valid  ,

            // manager 17, lane 18, stream 1      
            input   wire                                        std__mgr17__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane18_strm1_data        ,
            output  wire                                        mgr17__std__lane18_strm1_data_valid  ,

            // manager 17, lane 19, stream 0      
            input   wire                                        std__mgr17__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane19_strm0_data        ,
            output  wire                                        mgr17__std__lane19_strm0_data_valid  ,

            // manager 17, lane 19, stream 1      
            input   wire                                        std__mgr17__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane19_strm1_data        ,
            output  wire                                        mgr17__std__lane19_strm1_data_valid  ,

            // manager 17, lane 20, stream 0      
            input   wire                                        std__mgr17__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane20_strm0_data        ,
            output  wire                                        mgr17__std__lane20_strm0_data_valid  ,

            // manager 17, lane 20, stream 1      
            input   wire                                        std__mgr17__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane20_strm1_data        ,
            output  wire                                        mgr17__std__lane20_strm1_data_valid  ,

            // manager 17, lane 21, stream 0      
            input   wire                                        std__mgr17__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane21_strm0_data        ,
            output  wire                                        mgr17__std__lane21_strm0_data_valid  ,

            // manager 17, lane 21, stream 1      
            input   wire                                        std__mgr17__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane21_strm1_data        ,
            output  wire                                        mgr17__std__lane21_strm1_data_valid  ,

            // manager 17, lane 22, stream 0      
            input   wire                                        std__mgr17__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane22_strm0_data        ,
            output  wire                                        mgr17__std__lane22_strm0_data_valid  ,

            // manager 17, lane 22, stream 1      
            input   wire                                        std__mgr17__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane22_strm1_data        ,
            output  wire                                        mgr17__std__lane22_strm1_data_valid  ,

            // manager 17, lane 23, stream 0      
            input   wire                                        std__mgr17__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane23_strm0_data        ,
            output  wire                                        mgr17__std__lane23_strm0_data_valid  ,

            // manager 17, lane 23, stream 1      
            input   wire                                        std__mgr17__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane23_strm1_data        ,
            output  wire                                        mgr17__std__lane23_strm1_data_valid  ,

            // manager 17, lane 24, stream 0      
            input   wire                                        std__mgr17__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane24_strm0_data        ,
            output  wire                                        mgr17__std__lane24_strm0_data_valid  ,

            // manager 17, lane 24, stream 1      
            input   wire                                        std__mgr17__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane24_strm1_data        ,
            output  wire                                        mgr17__std__lane24_strm1_data_valid  ,

            // manager 17, lane 25, stream 0      
            input   wire                                        std__mgr17__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane25_strm0_data        ,
            output  wire                                        mgr17__std__lane25_strm0_data_valid  ,

            // manager 17, lane 25, stream 1      
            input   wire                                        std__mgr17__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane25_strm1_data        ,
            output  wire                                        mgr17__std__lane25_strm1_data_valid  ,

            // manager 17, lane 26, stream 0      
            input   wire                                        std__mgr17__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane26_strm0_data        ,
            output  wire                                        mgr17__std__lane26_strm0_data_valid  ,

            // manager 17, lane 26, stream 1      
            input   wire                                        std__mgr17__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane26_strm1_data        ,
            output  wire                                        mgr17__std__lane26_strm1_data_valid  ,

            // manager 17, lane 27, stream 0      
            input   wire                                        std__mgr17__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane27_strm0_data        ,
            output  wire                                        mgr17__std__lane27_strm0_data_valid  ,

            // manager 17, lane 27, stream 1      
            input   wire                                        std__mgr17__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane27_strm1_data        ,
            output  wire                                        mgr17__std__lane27_strm1_data_valid  ,

            // manager 17, lane 28, stream 0      
            input   wire                                        std__mgr17__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane28_strm0_data        ,
            output  wire                                        mgr17__std__lane28_strm0_data_valid  ,

            // manager 17, lane 28, stream 1      
            input   wire                                        std__mgr17__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane28_strm1_data        ,
            output  wire                                        mgr17__std__lane28_strm1_data_valid  ,

            // manager 17, lane 29, stream 0      
            input   wire                                        std__mgr17__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane29_strm0_data        ,
            output  wire                                        mgr17__std__lane29_strm0_data_valid  ,

            // manager 17, lane 29, stream 1      
            input   wire                                        std__mgr17__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane29_strm1_data        ,
            output  wire                                        mgr17__std__lane29_strm1_data_valid  ,

            // manager 17, lane 30, stream 0      
            input   wire                                        std__mgr17__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane30_strm0_data        ,
            output  wire                                        mgr17__std__lane30_strm0_data_valid  ,

            // manager 17, lane 30, stream 1      
            input   wire                                        std__mgr17__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane30_strm1_data        ,
            output  wire                                        mgr17__std__lane30_strm1_data_valid  ,

            // manager 17, lane 31, stream 0      
            input   wire                                        std__mgr17__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane31_strm0_data        ,
            output  wire                                        mgr17__std__lane31_strm0_data_valid  ,

            // manager 17, lane 31, stream 1      
            input   wire                                        std__mgr17__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr17__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr17__std__lane31_strm1_data        ,
            output  wire                                        mgr17__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 18, lane 0, stream 0      
            input   wire                                        std__mgr18__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane0_strm0_data        ,
            output  wire                                        mgr18__std__lane0_strm0_data_valid  ,

            // manager 18, lane 0, stream 1      
            input   wire                                        std__mgr18__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane0_strm1_data        ,
            output  wire                                        mgr18__std__lane0_strm1_data_valid  ,

            // manager 18, lane 1, stream 0      
            input   wire                                        std__mgr18__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane1_strm0_data        ,
            output  wire                                        mgr18__std__lane1_strm0_data_valid  ,

            // manager 18, lane 1, stream 1      
            input   wire                                        std__mgr18__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane1_strm1_data        ,
            output  wire                                        mgr18__std__lane1_strm1_data_valid  ,

            // manager 18, lane 2, stream 0      
            input   wire                                        std__mgr18__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane2_strm0_data        ,
            output  wire                                        mgr18__std__lane2_strm0_data_valid  ,

            // manager 18, lane 2, stream 1      
            input   wire                                        std__mgr18__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane2_strm1_data        ,
            output  wire                                        mgr18__std__lane2_strm1_data_valid  ,

            // manager 18, lane 3, stream 0      
            input   wire                                        std__mgr18__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane3_strm0_data        ,
            output  wire                                        mgr18__std__lane3_strm0_data_valid  ,

            // manager 18, lane 3, stream 1      
            input   wire                                        std__mgr18__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane3_strm1_data        ,
            output  wire                                        mgr18__std__lane3_strm1_data_valid  ,

            // manager 18, lane 4, stream 0      
            input   wire                                        std__mgr18__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane4_strm0_data        ,
            output  wire                                        mgr18__std__lane4_strm0_data_valid  ,

            // manager 18, lane 4, stream 1      
            input   wire                                        std__mgr18__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane4_strm1_data        ,
            output  wire                                        mgr18__std__lane4_strm1_data_valid  ,

            // manager 18, lane 5, stream 0      
            input   wire                                        std__mgr18__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane5_strm0_data        ,
            output  wire                                        mgr18__std__lane5_strm0_data_valid  ,

            // manager 18, lane 5, stream 1      
            input   wire                                        std__mgr18__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane5_strm1_data        ,
            output  wire                                        mgr18__std__lane5_strm1_data_valid  ,

            // manager 18, lane 6, stream 0      
            input   wire                                        std__mgr18__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane6_strm0_data        ,
            output  wire                                        mgr18__std__lane6_strm0_data_valid  ,

            // manager 18, lane 6, stream 1      
            input   wire                                        std__mgr18__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane6_strm1_data        ,
            output  wire                                        mgr18__std__lane6_strm1_data_valid  ,

            // manager 18, lane 7, stream 0      
            input   wire                                        std__mgr18__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane7_strm0_data        ,
            output  wire                                        mgr18__std__lane7_strm0_data_valid  ,

            // manager 18, lane 7, stream 1      
            input   wire                                        std__mgr18__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane7_strm1_data        ,
            output  wire                                        mgr18__std__lane7_strm1_data_valid  ,

            // manager 18, lane 8, stream 0      
            input   wire                                        std__mgr18__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane8_strm0_data        ,
            output  wire                                        mgr18__std__lane8_strm0_data_valid  ,

            // manager 18, lane 8, stream 1      
            input   wire                                        std__mgr18__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane8_strm1_data        ,
            output  wire                                        mgr18__std__lane8_strm1_data_valid  ,

            // manager 18, lane 9, stream 0      
            input   wire                                        std__mgr18__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane9_strm0_data        ,
            output  wire                                        mgr18__std__lane9_strm0_data_valid  ,

            // manager 18, lane 9, stream 1      
            input   wire                                        std__mgr18__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane9_strm1_data        ,
            output  wire                                        mgr18__std__lane9_strm1_data_valid  ,

            // manager 18, lane 10, stream 0      
            input   wire                                        std__mgr18__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane10_strm0_data        ,
            output  wire                                        mgr18__std__lane10_strm0_data_valid  ,

            // manager 18, lane 10, stream 1      
            input   wire                                        std__mgr18__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane10_strm1_data        ,
            output  wire                                        mgr18__std__lane10_strm1_data_valid  ,

            // manager 18, lane 11, stream 0      
            input   wire                                        std__mgr18__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane11_strm0_data        ,
            output  wire                                        mgr18__std__lane11_strm0_data_valid  ,

            // manager 18, lane 11, stream 1      
            input   wire                                        std__mgr18__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane11_strm1_data        ,
            output  wire                                        mgr18__std__lane11_strm1_data_valid  ,

            // manager 18, lane 12, stream 0      
            input   wire                                        std__mgr18__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane12_strm0_data        ,
            output  wire                                        mgr18__std__lane12_strm0_data_valid  ,

            // manager 18, lane 12, stream 1      
            input   wire                                        std__mgr18__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane12_strm1_data        ,
            output  wire                                        mgr18__std__lane12_strm1_data_valid  ,

            // manager 18, lane 13, stream 0      
            input   wire                                        std__mgr18__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane13_strm0_data        ,
            output  wire                                        mgr18__std__lane13_strm0_data_valid  ,

            // manager 18, lane 13, stream 1      
            input   wire                                        std__mgr18__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane13_strm1_data        ,
            output  wire                                        mgr18__std__lane13_strm1_data_valid  ,

            // manager 18, lane 14, stream 0      
            input   wire                                        std__mgr18__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane14_strm0_data        ,
            output  wire                                        mgr18__std__lane14_strm0_data_valid  ,

            // manager 18, lane 14, stream 1      
            input   wire                                        std__mgr18__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane14_strm1_data        ,
            output  wire                                        mgr18__std__lane14_strm1_data_valid  ,

            // manager 18, lane 15, stream 0      
            input   wire                                        std__mgr18__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane15_strm0_data        ,
            output  wire                                        mgr18__std__lane15_strm0_data_valid  ,

            // manager 18, lane 15, stream 1      
            input   wire                                        std__mgr18__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane15_strm1_data        ,
            output  wire                                        mgr18__std__lane15_strm1_data_valid  ,

            // manager 18, lane 16, stream 0      
            input   wire                                        std__mgr18__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane16_strm0_data        ,
            output  wire                                        mgr18__std__lane16_strm0_data_valid  ,

            // manager 18, lane 16, stream 1      
            input   wire                                        std__mgr18__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane16_strm1_data        ,
            output  wire                                        mgr18__std__lane16_strm1_data_valid  ,

            // manager 18, lane 17, stream 0      
            input   wire                                        std__mgr18__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane17_strm0_data        ,
            output  wire                                        mgr18__std__lane17_strm0_data_valid  ,

            // manager 18, lane 17, stream 1      
            input   wire                                        std__mgr18__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane17_strm1_data        ,
            output  wire                                        mgr18__std__lane17_strm1_data_valid  ,

            // manager 18, lane 18, stream 0      
            input   wire                                        std__mgr18__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane18_strm0_data        ,
            output  wire                                        mgr18__std__lane18_strm0_data_valid  ,

            // manager 18, lane 18, stream 1      
            input   wire                                        std__mgr18__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane18_strm1_data        ,
            output  wire                                        mgr18__std__lane18_strm1_data_valid  ,

            // manager 18, lane 19, stream 0      
            input   wire                                        std__mgr18__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane19_strm0_data        ,
            output  wire                                        mgr18__std__lane19_strm0_data_valid  ,

            // manager 18, lane 19, stream 1      
            input   wire                                        std__mgr18__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane19_strm1_data        ,
            output  wire                                        mgr18__std__lane19_strm1_data_valid  ,

            // manager 18, lane 20, stream 0      
            input   wire                                        std__mgr18__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane20_strm0_data        ,
            output  wire                                        mgr18__std__lane20_strm0_data_valid  ,

            // manager 18, lane 20, stream 1      
            input   wire                                        std__mgr18__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane20_strm1_data        ,
            output  wire                                        mgr18__std__lane20_strm1_data_valid  ,

            // manager 18, lane 21, stream 0      
            input   wire                                        std__mgr18__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane21_strm0_data        ,
            output  wire                                        mgr18__std__lane21_strm0_data_valid  ,

            // manager 18, lane 21, stream 1      
            input   wire                                        std__mgr18__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane21_strm1_data        ,
            output  wire                                        mgr18__std__lane21_strm1_data_valid  ,

            // manager 18, lane 22, stream 0      
            input   wire                                        std__mgr18__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane22_strm0_data        ,
            output  wire                                        mgr18__std__lane22_strm0_data_valid  ,

            // manager 18, lane 22, stream 1      
            input   wire                                        std__mgr18__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane22_strm1_data        ,
            output  wire                                        mgr18__std__lane22_strm1_data_valid  ,

            // manager 18, lane 23, stream 0      
            input   wire                                        std__mgr18__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane23_strm0_data        ,
            output  wire                                        mgr18__std__lane23_strm0_data_valid  ,

            // manager 18, lane 23, stream 1      
            input   wire                                        std__mgr18__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane23_strm1_data        ,
            output  wire                                        mgr18__std__lane23_strm1_data_valid  ,

            // manager 18, lane 24, stream 0      
            input   wire                                        std__mgr18__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane24_strm0_data        ,
            output  wire                                        mgr18__std__lane24_strm0_data_valid  ,

            // manager 18, lane 24, stream 1      
            input   wire                                        std__mgr18__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane24_strm1_data        ,
            output  wire                                        mgr18__std__lane24_strm1_data_valid  ,

            // manager 18, lane 25, stream 0      
            input   wire                                        std__mgr18__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane25_strm0_data        ,
            output  wire                                        mgr18__std__lane25_strm0_data_valid  ,

            // manager 18, lane 25, stream 1      
            input   wire                                        std__mgr18__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane25_strm1_data        ,
            output  wire                                        mgr18__std__lane25_strm1_data_valid  ,

            // manager 18, lane 26, stream 0      
            input   wire                                        std__mgr18__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane26_strm0_data        ,
            output  wire                                        mgr18__std__lane26_strm0_data_valid  ,

            // manager 18, lane 26, stream 1      
            input   wire                                        std__mgr18__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane26_strm1_data        ,
            output  wire                                        mgr18__std__lane26_strm1_data_valid  ,

            // manager 18, lane 27, stream 0      
            input   wire                                        std__mgr18__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane27_strm0_data        ,
            output  wire                                        mgr18__std__lane27_strm0_data_valid  ,

            // manager 18, lane 27, stream 1      
            input   wire                                        std__mgr18__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane27_strm1_data        ,
            output  wire                                        mgr18__std__lane27_strm1_data_valid  ,

            // manager 18, lane 28, stream 0      
            input   wire                                        std__mgr18__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane28_strm0_data        ,
            output  wire                                        mgr18__std__lane28_strm0_data_valid  ,

            // manager 18, lane 28, stream 1      
            input   wire                                        std__mgr18__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane28_strm1_data        ,
            output  wire                                        mgr18__std__lane28_strm1_data_valid  ,

            // manager 18, lane 29, stream 0      
            input   wire                                        std__mgr18__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane29_strm0_data        ,
            output  wire                                        mgr18__std__lane29_strm0_data_valid  ,

            // manager 18, lane 29, stream 1      
            input   wire                                        std__mgr18__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane29_strm1_data        ,
            output  wire                                        mgr18__std__lane29_strm1_data_valid  ,

            // manager 18, lane 30, stream 0      
            input   wire                                        std__mgr18__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane30_strm0_data        ,
            output  wire                                        mgr18__std__lane30_strm0_data_valid  ,

            // manager 18, lane 30, stream 1      
            input   wire                                        std__mgr18__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane30_strm1_data        ,
            output  wire                                        mgr18__std__lane30_strm1_data_valid  ,

            // manager 18, lane 31, stream 0      
            input   wire                                        std__mgr18__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane31_strm0_data        ,
            output  wire                                        mgr18__std__lane31_strm0_data_valid  ,

            // manager 18, lane 31, stream 1      
            input   wire                                        std__mgr18__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr18__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr18__std__lane31_strm1_data        ,
            output  wire                                        mgr18__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 19, lane 0, stream 0      
            input   wire                                        std__mgr19__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane0_strm0_data        ,
            output  wire                                        mgr19__std__lane0_strm0_data_valid  ,

            // manager 19, lane 0, stream 1      
            input   wire                                        std__mgr19__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane0_strm1_data        ,
            output  wire                                        mgr19__std__lane0_strm1_data_valid  ,

            // manager 19, lane 1, stream 0      
            input   wire                                        std__mgr19__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane1_strm0_data        ,
            output  wire                                        mgr19__std__lane1_strm0_data_valid  ,

            // manager 19, lane 1, stream 1      
            input   wire                                        std__mgr19__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane1_strm1_data        ,
            output  wire                                        mgr19__std__lane1_strm1_data_valid  ,

            // manager 19, lane 2, stream 0      
            input   wire                                        std__mgr19__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane2_strm0_data        ,
            output  wire                                        mgr19__std__lane2_strm0_data_valid  ,

            // manager 19, lane 2, stream 1      
            input   wire                                        std__mgr19__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane2_strm1_data        ,
            output  wire                                        mgr19__std__lane2_strm1_data_valid  ,

            // manager 19, lane 3, stream 0      
            input   wire                                        std__mgr19__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane3_strm0_data        ,
            output  wire                                        mgr19__std__lane3_strm0_data_valid  ,

            // manager 19, lane 3, stream 1      
            input   wire                                        std__mgr19__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane3_strm1_data        ,
            output  wire                                        mgr19__std__lane3_strm1_data_valid  ,

            // manager 19, lane 4, stream 0      
            input   wire                                        std__mgr19__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane4_strm0_data        ,
            output  wire                                        mgr19__std__lane4_strm0_data_valid  ,

            // manager 19, lane 4, stream 1      
            input   wire                                        std__mgr19__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane4_strm1_data        ,
            output  wire                                        mgr19__std__lane4_strm1_data_valid  ,

            // manager 19, lane 5, stream 0      
            input   wire                                        std__mgr19__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane5_strm0_data        ,
            output  wire                                        mgr19__std__lane5_strm0_data_valid  ,

            // manager 19, lane 5, stream 1      
            input   wire                                        std__mgr19__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane5_strm1_data        ,
            output  wire                                        mgr19__std__lane5_strm1_data_valid  ,

            // manager 19, lane 6, stream 0      
            input   wire                                        std__mgr19__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane6_strm0_data        ,
            output  wire                                        mgr19__std__lane6_strm0_data_valid  ,

            // manager 19, lane 6, stream 1      
            input   wire                                        std__mgr19__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane6_strm1_data        ,
            output  wire                                        mgr19__std__lane6_strm1_data_valid  ,

            // manager 19, lane 7, stream 0      
            input   wire                                        std__mgr19__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane7_strm0_data        ,
            output  wire                                        mgr19__std__lane7_strm0_data_valid  ,

            // manager 19, lane 7, stream 1      
            input   wire                                        std__mgr19__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane7_strm1_data        ,
            output  wire                                        mgr19__std__lane7_strm1_data_valid  ,

            // manager 19, lane 8, stream 0      
            input   wire                                        std__mgr19__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane8_strm0_data        ,
            output  wire                                        mgr19__std__lane8_strm0_data_valid  ,

            // manager 19, lane 8, stream 1      
            input   wire                                        std__mgr19__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane8_strm1_data        ,
            output  wire                                        mgr19__std__lane8_strm1_data_valid  ,

            // manager 19, lane 9, stream 0      
            input   wire                                        std__mgr19__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane9_strm0_data        ,
            output  wire                                        mgr19__std__lane9_strm0_data_valid  ,

            // manager 19, lane 9, stream 1      
            input   wire                                        std__mgr19__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane9_strm1_data        ,
            output  wire                                        mgr19__std__lane9_strm1_data_valid  ,

            // manager 19, lane 10, stream 0      
            input   wire                                        std__mgr19__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane10_strm0_data        ,
            output  wire                                        mgr19__std__lane10_strm0_data_valid  ,

            // manager 19, lane 10, stream 1      
            input   wire                                        std__mgr19__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane10_strm1_data        ,
            output  wire                                        mgr19__std__lane10_strm1_data_valid  ,

            // manager 19, lane 11, stream 0      
            input   wire                                        std__mgr19__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane11_strm0_data        ,
            output  wire                                        mgr19__std__lane11_strm0_data_valid  ,

            // manager 19, lane 11, stream 1      
            input   wire                                        std__mgr19__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane11_strm1_data        ,
            output  wire                                        mgr19__std__lane11_strm1_data_valid  ,

            // manager 19, lane 12, stream 0      
            input   wire                                        std__mgr19__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane12_strm0_data        ,
            output  wire                                        mgr19__std__lane12_strm0_data_valid  ,

            // manager 19, lane 12, stream 1      
            input   wire                                        std__mgr19__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane12_strm1_data        ,
            output  wire                                        mgr19__std__lane12_strm1_data_valid  ,

            // manager 19, lane 13, stream 0      
            input   wire                                        std__mgr19__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane13_strm0_data        ,
            output  wire                                        mgr19__std__lane13_strm0_data_valid  ,

            // manager 19, lane 13, stream 1      
            input   wire                                        std__mgr19__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane13_strm1_data        ,
            output  wire                                        mgr19__std__lane13_strm1_data_valid  ,

            // manager 19, lane 14, stream 0      
            input   wire                                        std__mgr19__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane14_strm0_data        ,
            output  wire                                        mgr19__std__lane14_strm0_data_valid  ,

            // manager 19, lane 14, stream 1      
            input   wire                                        std__mgr19__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane14_strm1_data        ,
            output  wire                                        mgr19__std__lane14_strm1_data_valid  ,

            // manager 19, lane 15, stream 0      
            input   wire                                        std__mgr19__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane15_strm0_data        ,
            output  wire                                        mgr19__std__lane15_strm0_data_valid  ,

            // manager 19, lane 15, stream 1      
            input   wire                                        std__mgr19__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane15_strm1_data        ,
            output  wire                                        mgr19__std__lane15_strm1_data_valid  ,

            // manager 19, lane 16, stream 0      
            input   wire                                        std__mgr19__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane16_strm0_data        ,
            output  wire                                        mgr19__std__lane16_strm0_data_valid  ,

            // manager 19, lane 16, stream 1      
            input   wire                                        std__mgr19__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane16_strm1_data        ,
            output  wire                                        mgr19__std__lane16_strm1_data_valid  ,

            // manager 19, lane 17, stream 0      
            input   wire                                        std__mgr19__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane17_strm0_data        ,
            output  wire                                        mgr19__std__lane17_strm0_data_valid  ,

            // manager 19, lane 17, stream 1      
            input   wire                                        std__mgr19__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane17_strm1_data        ,
            output  wire                                        mgr19__std__lane17_strm1_data_valid  ,

            // manager 19, lane 18, stream 0      
            input   wire                                        std__mgr19__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane18_strm0_data        ,
            output  wire                                        mgr19__std__lane18_strm0_data_valid  ,

            // manager 19, lane 18, stream 1      
            input   wire                                        std__mgr19__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane18_strm1_data        ,
            output  wire                                        mgr19__std__lane18_strm1_data_valid  ,

            // manager 19, lane 19, stream 0      
            input   wire                                        std__mgr19__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane19_strm0_data        ,
            output  wire                                        mgr19__std__lane19_strm0_data_valid  ,

            // manager 19, lane 19, stream 1      
            input   wire                                        std__mgr19__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane19_strm1_data        ,
            output  wire                                        mgr19__std__lane19_strm1_data_valid  ,

            // manager 19, lane 20, stream 0      
            input   wire                                        std__mgr19__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane20_strm0_data        ,
            output  wire                                        mgr19__std__lane20_strm0_data_valid  ,

            // manager 19, lane 20, stream 1      
            input   wire                                        std__mgr19__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane20_strm1_data        ,
            output  wire                                        mgr19__std__lane20_strm1_data_valid  ,

            // manager 19, lane 21, stream 0      
            input   wire                                        std__mgr19__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane21_strm0_data        ,
            output  wire                                        mgr19__std__lane21_strm0_data_valid  ,

            // manager 19, lane 21, stream 1      
            input   wire                                        std__mgr19__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane21_strm1_data        ,
            output  wire                                        mgr19__std__lane21_strm1_data_valid  ,

            // manager 19, lane 22, stream 0      
            input   wire                                        std__mgr19__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane22_strm0_data        ,
            output  wire                                        mgr19__std__lane22_strm0_data_valid  ,

            // manager 19, lane 22, stream 1      
            input   wire                                        std__mgr19__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane22_strm1_data        ,
            output  wire                                        mgr19__std__lane22_strm1_data_valid  ,

            // manager 19, lane 23, stream 0      
            input   wire                                        std__mgr19__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane23_strm0_data        ,
            output  wire                                        mgr19__std__lane23_strm0_data_valid  ,

            // manager 19, lane 23, stream 1      
            input   wire                                        std__mgr19__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane23_strm1_data        ,
            output  wire                                        mgr19__std__lane23_strm1_data_valid  ,

            // manager 19, lane 24, stream 0      
            input   wire                                        std__mgr19__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane24_strm0_data        ,
            output  wire                                        mgr19__std__lane24_strm0_data_valid  ,

            // manager 19, lane 24, stream 1      
            input   wire                                        std__mgr19__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane24_strm1_data        ,
            output  wire                                        mgr19__std__lane24_strm1_data_valid  ,

            // manager 19, lane 25, stream 0      
            input   wire                                        std__mgr19__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane25_strm0_data        ,
            output  wire                                        mgr19__std__lane25_strm0_data_valid  ,

            // manager 19, lane 25, stream 1      
            input   wire                                        std__mgr19__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane25_strm1_data        ,
            output  wire                                        mgr19__std__lane25_strm1_data_valid  ,

            // manager 19, lane 26, stream 0      
            input   wire                                        std__mgr19__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane26_strm0_data        ,
            output  wire                                        mgr19__std__lane26_strm0_data_valid  ,

            // manager 19, lane 26, stream 1      
            input   wire                                        std__mgr19__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane26_strm1_data        ,
            output  wire                                        mgr19__std__lane26_strm1_data_valid  ,

            // manager 19, lane 27, stream 0      
            input   wire                                        std__mgr19__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane27_strm0_data        ,
            output  wire                                        mgr19__std__lane27_strm0_data_valid  ,

            // manager 19, lane 27, stream 1      
            input   wire                                        std__mgr19__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane27_strm1_data        ,
            output  wire                                        mgr19__std__lane27_strm1_data_valid  ,

            // manager 19, lane 28, stream 0      
            input   wire                                        std__mgr19__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane28_strm0_data        ,
            output  wire                                        mgr19__std__lane28_strm0_data_valid  ,

            // manager 19, lane 28, stream 1      
            input   wire                                        std__mgr19__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane28_strm1_data        ,
            output  wire                                        mgr19__std__lane28_strm1_data_valid  ,

            // manager 19, lane 29, stream 0      
            input   wire                                        std__mgr19__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane29_strm0_data        ,
            output  wire                                        mgr19__std__lane29_strm0_data_valid  ,

            // manager 19, lane 29, stream 1      
            input   wire                                        std__mgr19__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane29_strm1_data        ,
            output  wire                                        mgr19__std__lane29_strm1_data_valid  ,

            // manager 19, lane 30, stream 0      
            input   wire                                        std__mgr19__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane30_strm0_data        ,
            output  wire                                        mgr19__std__lane30_strm0_data_valid  ,

            // manager 19, lane 30, stream 1      
            input   wire                                        std__mgr19__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane30_strm1_data        ,
            output  wire                                        mgr19__std__lane30_strm1_data_valid  ,

            // manager 19, lane 31, stream 0      
            input   wire                                        std__mgr19__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane31_strm0_data        ,
            output  wire                                        mgr19__std__lane31_strm0_data_valid  ,

            // manager 19, lane 31, stream 1      
            input   wire                                        std__mgr19__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr19__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr19__std__lane31_strm1_data        ,
            output  wire                                        mgr19__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 20, lane 0, stream 0      
            input   wire                                        std__mgr20__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane0_strm0_data        ,
            output  wire                                        mgr20__std__lane0_strm0_data_valid  ,

            // manager 20, lane 0, stream 1      
            input   wire                                        std__mgr20__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane0_strm1_data        ,
            output  wire                                        mgr20__std__lane0_strm1_data_valid  ,

            // manager 20, lane 1, stream 0      
            input   wire                                        std__mgr20__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane1_strm0_data        ,
            output  wire                                        mgr20__std__lane1_strm0_data_valid  ,

            // manager 20, lane 1, stream 1      
            input   wire                                        std__mgr20__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane1_strm1_data        ,
            output  wire                                        mgr20__std__lane1_strm1_data_valid  ,

            // manager 20, lane 2, stream 0      
            input   wire                                        std__mgr20__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane2_strm0_data        ,
            output  wire                                        mgr20__std__lane2_strm0_data_valid  ,

            // manager 20, lane 2, stream 1      
            input   wire                                        std__mgr20__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane2_strm1_data        ,
            output  wire                                        mgr20__std__lane2_strm1_data_valid  ,

            // manager 20, lane 3, stream 0      
            input   wire                                        std__mgr20__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane3_strm0_data        ,
            output  wire                                        mgr20__std__lane3_strm0_data_valid  ,

            // manager 20, lane 3, stream 1      
            input   wire                                        std__mgr20__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane3_strm1_data        ,
            output  wire                                        mgr20__std__lane3_strm1_data_valid  ,

            // manager 20, lane 4, stream 0      
            input   wire                                        std__mgr20__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane4_strm0_data        ,
            output  wire                                        mgr20__std__lane4_strm0_data_valid  ,

            // manager 20, lane 4, stream 1      
            input   wire                                        std__mgr20__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane4_strm1_data        ,
            output  wire                                        mgr20__std__lane4_strm1_data_valid  ,

            // manager 20, lane 5, stream 0      
            input   wire                                        std__mgr20__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane5_strm0_data        ,
            output  wire                                        mgr20__std__lane5_strm0_data_valid  ,

            // manager 20, lane 5, stream 1      
            input   wire                                        std__mgr20__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane5_strm1_data        ,
            output  wire                                        mgr20__std__lane5_strm1_data_valid  ,

            // manager 20, lane 6, stream 0      
            input   wire                                        std__mgr20__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane6_strm0_data        ,
            output  wire                                        mgr20__std__lane6_strm0_data_valid  ,

            // manager 20, lane 6, stream 1      
            input   wire                                        std__mgr20__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane6_strm1_data        ,
            output  wire                                        mgr20__std__lane6_strm1_data_valid  ,

            // manager 20, lane 7, stream 0      
            input   wire                                        std__mgr20__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane7_strm0_data        ,
            output  wire                                        mgr20__std__lane7_strm0_data_valid  ,

            // manager 20, lane 7, stream 1      
            input   wire                                        std__mgr20__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane7_strm1_data        ,
            output  wire                                        mgr20__std__lane7_strm1_data_valid  ,

            // manager 20, lane 8, stream 0      
            input   wire                                        std__mgr20__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane8_strm0_data        ,
            output  wire                                        mgr20__std__lane8_strm0_data_valid  ,

            // manager 20, lane 8, stream 1      
            input   wire                                        std__mgr20__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane8_strm1_data        ,
            output  wire                                        mgr20__std__lane8_strm1_data_valid  ,

            // manager 20, lane 9, stream 0      
            input   wire                                        std__mgr20__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane9_strm0_data        ,
            output  wire                                        mgr20__std__lane9_strm0_data_valid  ,

            // manager 20, lane 9, stream 1      
            input   wire                                        std__mgr20__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane9_strm1_data        ,
            output  wire                                        mgr20__std__lane9_strm1_data_valid  ,

            // manager 20, lane 10, stream 0      
            input   wire                                        std__mgr20__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane10_strm0_data        ,
            output  wire                                        mgr20__std__lane10_strm0_data_valid  ,

            // manager 20, lane 10, stream 1      
            input   wire                                        std__mgr20__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane10_strm1_data        ,
            output  wire                                        mgr20__std__lane10_strm1_data_valid  ,

            // manager 20, lane 11, stream 0      
            input   wire                                        std__mgr20__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane11_strm0_data        ,
            output  wire                                        mgr20__std__lane11_strm0_data_valid  ,

            // manager 20, lane 11, stream 1      
            input   wire                                        std__mgr20__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane11_strm1_data        ,
            output  wire                                        mgr20__std__lane11_strm1_data_valid  ,

            // manager 20, lane 12, stream 0      
            input   wire                                        std__mgr20__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane12_strm0_data        ,
            output  wire                                        mgr20__std__lane12_strm0_data_valid  ,

            // manager 20, lane 12, stream 1      
            input   wire                                        std__mgr20__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane12_strm1_data        ,
            output  wire                                        mgr20__std__lane12_strm1_data_valid  ,

            // manager 20, lane 13, stream 0      
            input   wire                                        std__mgr20__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane13_strm0_data        ,
            output  wire                                        mgr20__std__lane13_strm0_data_valid  ,

            // manager 20, lane 13, stream 1      
            input   wire                                        std__mgr20__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane13_strm1_data        ,
            output  wire                                        mgr20__std__lane13_strm1_data_valid  ,

            // manager 20, lane 14, stream 0      
            input   wire                                        std__mgr20__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane14_strm0_data        ,
            output  wire                                        mgr20__std__lane14_strm0_data_valid  ,

            // manager 20, lane 14, stream 1      
            input   wire                                        std__mgr20__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane14_strm1_data        ,
            output  wire                                        mgr20__std__lane14_strm1_data_valid  ,

            // manager 20, lane 15, stream 0      
            input   wire                                        std__mgr20__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane15_strm0_data        ,
            output  wire                                        mgr20__std__lane15_strm0_data_valid  ,

            // manager 20, lane 15, stream 1      
            input   wire                                        std__mgr20__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane15_strm1_data        ,
            output  wire                                        mgr20__std__lane15_strm1_data_valid  ,

            // manager 20, lane 16, stream 0      
            input   wire                                        std__mgr20__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane16_strm0_data        ,
            output  wire                                        mgr20__std__lane16_strm0_data_valid  ,

            // manager 20, lane 16, stream 1      
            input   wire                                        std__mgr20__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane16_strm1_data        ,
            output  wire                                        mgr20__std__lane16_strm1_data_valid  ,

            // manager 20, lane 17, stream 0      
            input   wire                                        std__mgr20__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane17_strm0_data        ,
            output  wire                                        mgr20__std__lane17_strm0_data_valid  ,

            // manager 20, lane 17, stream 1      
            input   wire                                        std__mgr20__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane17_strm1_data        ,
            output  wire                                        mgr20__std__lane17_strm1_data_valid  ,

            // manager 20, lane 18, stream 0      
            input   wire                                        std__mgr20__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane18_strm0_data        ,
            output  wire                                        mgr20__std__lane18_strm0_data_valid  ,

            // manager 20, lane 18, stream 1      
            input   wire                                        std__mgr20__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane18_strm1_data        ,
            output  wire                                        mgr20__std__lane18_strm1_data_valid  ,

            // manager 20, lane 19, stream 0      
            input   wire                                        std__mgr20__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane19_strm0_data        ,
            output  wire                                        mgr20__std__lane19_strm0_data_valid  ,

            // manager 20, lane 19, stream 1      
            input   wire                                        std__mgr20__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane19_strm1_data        ,
            output  wire                                        mgr20__std__lane19_strm1_data_valid  ,

            // manager 20, lane 20, stream 0      
            input   wire                                        std__mgr20__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane20_strm0_data        ,
            output  wire                                        mgr20__std__lane20_strm0_data_valid  ,

            // manager 20, lane 20, stream 1      
            input   wire                                        std__mgr20__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane20_strm1_data        ,
            output  wire                                        mgr20__std__lane20_strm1_data_valid  ,

            // manager 20, lane 21, stream 0      
            input   wire                                        std__mgr20__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane21_strm0_data        ,
            output  wire                                        mgr20__std__lane21_strm0_data_valid  ,

            // manager 20, lane 21, stream 1      
            input   wire                                        std__mgr20__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane21_strm1_data        ,
            output  wire                                        mgr20__std__lane21_strm1_data_valid  ,

            // manager 20, lane 22, stream 0      
            input   wire                                        std__mgr20__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane22_strm0_data        ,
            output  wire                                        mgr20__std__lane22_strm0_data_valid  ,

            // manager 20, lane 22, stream 1      
            input   wire                                        std__mgr20__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane22_strm1_data        ,
            output  wire                                        mgr20__std__lane22_strm1_data_valid  ,

            // manager 20, lane 23, stream 0      
            input   wire                                        std__mgr20__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane23_strm0_data        ,
            output  wire                                        mgr20__std__lane23_strm0_data_valid  ,

            // manager 20, lane 23, stream 1      
            input   wire                                        std__mgr20__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane23_strm1_data        ,
            output  wire                                        mgr20__std__lane23_strm1_data_valid  ,

            // manager 20, lane 24, stream 0      
            input   wire                                        std__mgr20__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane24_strm0_data        ,
            output  wire                                        mgr20__std__lane24_strm0_data_valid  ,

            // manager 20, lane 24, stream 1      
            input   wire                                        std__mgr20__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane24_strm1_data        ,
            output  wire                                        mgr20__std__lane24_strm1_data_valid  ,

            // manager 20, lane 25, stream 0      
            input   wire                                        std__mgr20__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane25_strm0_data        ,
            output  wire                                        mgr20__std__lane25_strm0_data_valid  ,

            // manager 20, lane 25, stream 1      
            input   wire                                        std__mgr20__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane25_strm1_data        ,
            output  wire                                        mgr20__std__lane25_strm1_data_valid  ,

            // manager 20, lane 26, stream 0      
            input   wire                                        std__mgr20__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane26_strm0_data        ,
            output  wire                                        mgr20__std__lane26_strm0_data_valid  ,

            // manager 20, lane 26, stream 1      
            input   wire                                        std__mgr20__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane26_strm1_data        ,
            output  wire                                        mgr20__std__lane26_strm1_data_valid  ,

            // manager 20, lane 27, stream 0      
            input   wire                                        std__mgr20__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane27_strm0_data        ,
            output  wire                                        mgr20__std__lane27_strm0_data_valid  ,

            // manager 20, lane 27, stream 1      
            input   wire                                        std__mgr20__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane27_strm1_data        ,
            output  wire                                        mgr20__std__lane27_strm1_data_valid  ,

            // manager 20, lane 28, stream 0      
            input   wire                                        std__mgr20__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane28_strm0_data        ,
            output  wire                                        mgr20__std__lane28_strm0_data_valid  ,

            // manager 20, lane 28, stream 1      
            input   wire                                        std__mgr20__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane28_strm1_data        ,
            output  wire                                        mgr20__std__lane28_strm1_data_valid  ,

            // manager 20, lane 29, stream 0      
            input   wire                                        std__mgr20__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane29_strm0_data        ,
            output  wire                                        mgr20__std__lane29_strm0_data_valid  ,

            // manager 20, lane 29, stream 1      
            input   wire                                        std__mgr20__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane29_strm1_data        ,
            output  wire                                        mgr20__std__lane29_strm1_data_valid  ,

            // manager 20, lane 30, stream 0      
            input   wire                                        std__mgr20__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane30_strm0_data        ,
            output  wire                                        mgr20__std__lane30_strm0_data_valid  ,

            // manager 20, lane 30, stream 1      
            input   wire                                        std__mgr20__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane30_strm1_data        ,
            output  wire                                        mgr20__std__lane30_strm1_data_valid  ,

            // manager 20, lane 31, stream 0      
            input   wire                                        std__mgr20__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane31_strm0_data        ,
            output  wire                                        mgr20__std__lane31_strm0_data_valid  ,

            // manager 20, lane 31, stream 1      
            input   wire                                        std__mgr20__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr20__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr20__std__lane31_strm1_data        ,
            output  wire                                        mgr20__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 21, lane 0, stream 0      
            input   wire                                        std__mgr21__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane0_strm0_data        ,
            output  wire                                        mgr21__std__lane0_strm0_data_valid  ,

            // manager 21, lane 0, stream 1      
            input   wire                                        std__mgr21__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane0_strm1_data        ,
            output  wire                                        mgr21__std__lane0_strm1_data_valid  ,

            // manager 21, lane 1, stream 0      
            input   wire                                        std__mgr21__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane1_strm0_data        ,
            output  wire                                        mgr21__std__lane1_strm0_data_valid  ,

            // manager 21, lane 1, stream 1      
            input   wire                                        std__mgr21__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane1_strm1_data        ,
            output  wire                                        mgr21__std__lane1_strm1_data_valid  ,

            // manager 21, lane 2, stream 0      
            input   wire                                        std__mgr21__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane2_strm0_data        ,
            output  wire                                        mgr21__std__lane2_strm0_data_valid  ,

            // manager 21, lane 2, stream 1      
            input   wire                                        std__mgr21__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane2_strm1_data        ,
            output  wire                                        mgr21__std__lane2_strm1_data_valid  ,

            // manager 21, lane 3, stream 0      
            input   wire                                        std__mgr21__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane3_strm0_data        ,
            output  wire                                        mgr21__std__lane3_strm0_data_valid  ,

            // manager 21, lane 3, stream 1      
            input   wire                                        std__mgr21__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane3_strm1_data        ,
            output  wire                                        mgr21__std__lane3_strm1_data_valid  ,

            // manager 21, lane 4, stream 0      
            input   wire                                        std__mgr21__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane4_strm0_data        ,
            output  wire                                        mgr21__std__lane4_strm0_data_valid  ,

            // manager 21, lane 4, stream 1      
            input   wire                                        std__mgr21__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane4_strm1_data        ,
            output  wire                                        mgr21__std__lane4_strm1_data_valid  ,

            // manager 21, lane 5, stream 0      
            input   wire                                        std__mgr21__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane5_strm0_data        ,
            output  wire                                        mgr21__std__lane5_strm0_data_valid  ,

            // manager 21, lane 5, stream 1      
            input   wire                                        std__mgr21__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane5_strm1_data        ,
            output  wire                                        mgr21__std__lane5_strm1_data_valid  ,

            // manager 21, lane 6, stream 0      
            input   wire                                        std__mgr21__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane6_strm0_data        ,
            output  wire                                        mgr21__std__lane6_strm0_data_valid  ,

            // manager 21, lane 6, stream 1      
            input   wire                                        std__mgr21__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane6_strm1_data        ,
            output  wire                                        mgr21__std__lane6_strm1_data_valid  ,

            // manager 21, lane 7, stream 0      
            input   wire                                        std__mgr21__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane7_strm0_data        ,
            output  wire                                        mgr21__std__lane7_strm0_data_valid  ,

            // manager 21, lane 7, stream 1      
            input   wire                                        std__mgr21__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane7_strm1_data        ,
            output  wire                                        mgr21__std__lane7_strm1_data_valid  ,

            // manager 21, lane 8, stream 0      
            input   wire                                        std__mgr21__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane8_strm0_data        ,
            output  wire                                        mgr21__std__lane8_strm0_data_valid  ,

            // manager 21, lane 8, stream 1      
            input   wire                                        std__mgr21__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane8_strm1_data        ,
            output  wire                                        mgr21__std__lane8_strm1_data_valid  ,

            // manager 21, lane 9, stream 0      
            input   wire                                        std__mgr21__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane9_strm0_data        ,
            output  wire                                        mgr21__std__lane9_strm0_data_valid  ,

            // manager 21, lane 9, stream 1      
            input   wire                                        std__mgr21__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane9_strm1_data        ,
            output  wire                                        mgr21__std__lane9_strm1_data_valid  ,

            // manager 21, lane 10, stream 0      
            input   wire                                        std__mgr21__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane10_strm0_data        ,
            output  wire                                        mgr21__std__lane10_strm0_data_valid  ,

            // manager 21, lane 10, stream 1      
            input   wire                                        std__mgr21__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane10_strm1_data        ,
            output  wire                                        mgr21__std__lane10_strm1_data_valid  ,

            // manager 21, lane 11, stream 0      
            input   wire                                        std__mgr21__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane11_strm0_data        ,
            output  wire                                        mgr21__std__lane11_strm0_data_valid  ,

            // manager 21, lane 11, stream 1      
            input   wire                                        std__mgr21__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane11_strm1_data        ,
            output  wire                                        mgr21__std__lane11_strm1_data_valid  ,

            // manager 21, lane 12, stream 0      
            input   wire                                        std__mgr21__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane12_strm0_data        ,
            output  wire                                        mgr21__std__lane12_strm0_data_valid  ,

            // manager 21, lane 12, stream 1      
            input   wire                                        std__mgr21__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane12_strm1_data        ,
            output  wire                                        mgr21__std__lane12_strm1_data_valid  ,

            // manager 21, lane 13, stream 0      
            input   wire                                        std__mgr21__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane13_strm0_data        ,
            output  wire                                        mgr21__std__lane13_strm0_data_valid  ,

            // manager 21, lane 13, stream 1      
            input   wire                                        std__mgr21__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane13_strm1_data        ,
            output  wire                                        mgr21__std__lane13_strm1_data_valid  ,

            // manager 21, lane 14, stream 0      
            input   wire                                        std__mgr21__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane14_strm0_data        ,
            output  wire                                        mgr21__std__lane14_strm0_data_valid  ,

            // manager 21, lane 14, stream 1      
            input   wire                                        std__mgr21__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane14_strm1_data        ,
            output  wire                                        mgr21__std__lane14_strm1_data_valid  ,

            // manager 21, lane 15, stream 0      
            input   wire                                        std__mgr21__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane15_strm0_data        ,
            output  wire                                        mgr21__std__lane15_strm0_data_valid  ,

            // manager 21, lane 15, stream 1      
            input   wire                                        std__mgr21__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane15_strm1_data        ,
            output  wire                                        mgr21__std__lane15_strm1_data_valid  ,

            // manager 21, lane 16, stream 0      
            input   wire                                        std__mgr21__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane16_strm0_data        ,
            output  wire                                        mgr21__std__lane16_strm0_data_valid  ,

            // manager 21, lane 16, stream 1      
            input   wire                                        std__mgr21__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane16_strm1_data        ,
            output  wire                                        mgr21__std__lane16_strm1_data_valid  ,

            // manager 21, lane 17, stream 0      
            input   wire                                        std__mgr21__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane17_strm0_data        ,
            output  wire                                        mgr21__std__lane17_strm0_data_valid  ,

            // manager 21, lane 17, stream 1      
            input   wire                                        std__mgr21__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane17_strm1_data        ,
            output  wire                                        mgr21__std__lane17_strm1_data_valid  ,

            // manager 21, lane 18, stream 0      
            input   wire                                        std__mgr21__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane18_strm0_data        ,
            output  wire                                        mgr21__std__lane18_strm0_data_valid  ,

            // manager 21, lane 18, stream 1      
            input   wire                                        std__mgr21__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane18_strm1_data        ,
            output  wire                                        mgr21__std__lane18_strm1_data_valid  ,

            // manager 21, lane 19, stream 0      
            input   wire                                        std__mgr21__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane19_strm0_data        ,
            output  wire                                        mgr21__std__lane19_strm0_data_valid  ,

            // manager 21, lane 19, stream 1      
            input   wire                                        std__mgr21__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane19_strm1_data        ,
            output  wire                                        mgr21__std__lane19_strm1_data_valid  ,

            // manager 21, lane 20, stream 0      
            input   wire                                        std__mgr21__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane20_strm0_data        ,
            output  wire                                        mgr21__std__lane20_strm0_data_valid  ,

            // manager 21, lane 20, stream 1      
            input   wire                                        std__mgr21__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane20_strm1_data        ,
            output  wire                                        mgr21__std__lane20_strm1_data_valid  ,

            // manager 21, lane 21, stream 0      
            input   wire                                        std__mgr21__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane21_strm0_data        ,
            output  wire                                        mgr21__std__lane21_strm0_data_valid  ,

            // manager 21, lane 21, stream 1      
            input   wire                                        std__mgr21__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane21_strm1_data        ,
            output  wire                                        mgr21__std__lane21_strm1_data_valid  ,

            // manager 21, lane 22, stream 0      
            input   wire                                        std__mgr21__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane22_strm0_data        ,
            output  wire                                        mgr21__std__lane22_strm0_data_valid  ,

            // manager 21, lane 22, stream 1      
            input   wire                                        std__mgr21__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane22_strm1_data        ,
            output  wire                                        mgr21__std__lane22_strm1_data_valid  ,

            // manager 21, lane 23, stream 0      
            input   wire                                        std__mgr21__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane23_strm0_data        ,
            output  wire                                        mgr21__std__lane23_strm0_data_valid  ,

            // manager 21, lane 23, stream 1      
            input   wire                                        std__mgr21__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane23_strm1_data        ,
            output  wire                                        mgr21__std__lane23_strm1_data_valid  ,

            // manager 21, lane 24, stream 0      
            input   wire                                        std__mgr21__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane24_strm0_data        ,
            output  wire                                        mgr21__std__lane24_strm0_data_valid  ,

            // manager 21, lane 24, stream 1      
            input   wire                                        std__mgr21__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane24_strm1_data        ,
            output  wire                                        mgr21__std__lane24_strm1_data_valid  ,

            // manager 21, lane 25, stream 0      
            input   wire                                        std__mgr21__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane25_strm0_data        ,
            output  wire                                        mgr21__std__lane25_strm0_data_valid  ,

            // manager 21, lane 25, stream 1      
            input   wire                                        std__mgr21__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane25_strm1_data        ,
            output  wire                                        mgr21__std__lane25_strm1_data_valid  ,

            // manager 21, lane 26, stream 0      
            input   wire                                        std__mgr21__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane26_strm0_data        ,
            output  wire                                        mgr21__std__lane26_strm0_data_valid  ,

            // manager 21, lane 26, stream 1      
            input   wire                                        std__mgr21__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane26_strm1_data        ,
            output  wire                                        mgr21__std__lane26_strm1_data_valid  ,

            // manager 21, lane 27, stream 0      
            input   wire                                        std__mgr21__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane27_strm0_data        ,
            output  wire                                        mgr21__std__lane27_strm0_data_valid  ,

            // manager 21, lane 27, stream 1      
            input   wire                                        std__mgr21__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane27_strm1_data        ,
            output  wire                                        mgr21__std__lane27_strm1_data_valid  ,

            // manager 21, lane 28, stream 0      
            input   wire                                        std__mgr21__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane28_strm0_data        ,
            output  wire                                        mgr21__std__lane28_strm0_data_valid  ,

            // manager 21, lane 28, stream 1      
            input   wire                                        std__mgr21__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane28_strm1_data        ,
            output  wire                                        mgr21__std__lane28_strm1_data_valid  ,

            // manager 21, lane 29, stream 0      
            input   wire                                        std__mgr21__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane29_strm0_data        ,
            output  wire                                        mgr21__std__lane29_strm0_data_valid  ,

            // manager 21, lane 29, stream 1      
            input   wire                                        std__mgr21__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane29_strm1_data        ,
            output  wire                                        mgr21__std__lane29_strm1_data_valid  ,

            // manager 21, lane 30, stream 0      
            input   wire                                        std__mgr21__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane30_strm0_data        ,
            output  wire                                        mgr21__std__lane30_strm0_data_valid  ,

            // manager 21, lane 30, stream 1      
            input   wire                                        std__mgr21__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane30_strm1_data        ,
            output  wire                                        mgr21__std__lane30_strm1_data_valid  ,

            // manager 21, lane 31, stream 0      
            input   wire                                        std__mgr21__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane31_strm0_data        ,
            output  wire                                        mgr21__std__lane31_strm0_data_valid  ,

            // manager 21, lane 31, stream 1      
            input   wire                                        std__mgr21__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr21__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr21__std__lane31_strm1_data        ,
            output  wire                                        mgr21__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 22, lane 0, stream 0      
            input   wire                                        std__mgr22__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane0_strm0_data        ,
            output  wire                                        mgr22__std__lane0_strm0_data_valid  ,

            // manager 22, lane 0, stream 1      
            input   wire                                        std__mgr22__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane0_strm1_data        ,
            output  wire                                        mgr22__std__lane0_strm1_data_valid  ,

            // manager 22, lane 1, stream 0      
            input   wire                                        std__mgr22__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane1_strm0_data        ,
            output  wire                                        mgr22__std__lane1_strm0_data_valid  ,

            // manager 22, lane 1, stream 1      
            input   wire                                        std__mgr22__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane1_strm1_data        ,
            output  wire                                        mgr22__std__lane1_strm1_data_valid  ,

            // manager 22, lane 2, stream 0      
            input   wire                                        std__mgr22__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane2_strm0_data        ,
            output  wire                                        mgr22__std__lane2_strm0_data_valid  ,

            // manager 22, lane 2, stream 1      
            input   wire                                        std__mgr22__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane2_strm1_data        ,
            output  wire                                        mgr22__std__lane2_strm1_data_valid  ,

            // manager 22, lane 3, stream 0      
            input   wire                                        std__mgr22__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane3_strm0_data        ,
            output  wire                                        mgr22__std__lane3_strm0_data_valid  ,

            // manager 22, lane 3, stream 1      
            input   wire                                        std__mgr22__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane3_strm1_data        ,
            output  wire                                        mgr22__std__lane3_strm1_data_valid  ,

            // manager 22, lane 4, stream 0      
            input   wire                                        std__mgr22__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane4_strm0_data        ,
            output  wire                                        mgr22__std__lane4_strm0_data_valid  ,

            // manager 22, lane 4, stream 1      
            input   wire                                        std__mgr22__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane4_strm1_data        ,
            output  wire                                        mgr22__std__lane4_strm1_data_valid  ,

            // manager 22, lane 5, stream 0      
            input   wire                                        std__mgr22__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane5_strm0_data        ,
            output  wire                                        mgr22__std__lane5_strm0_data_valid  ,

            // manager 22, lane 5, stream 1      
            input   wire                                        std__mgr22__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane5_strm1_data        ,
            output  wire                                        mgr22__std__lane5_strm1_data_valid  ,

            // manager 22, lane 6, stream 0      
            input   wire                                        std__mgr22__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane6_strm0_data        ,
            output  wire                                        mgr22__std__lane6_strm0_data_valid  ,

            // manager 22, lane 6, stream 1      
            input   wire                                        std__mgr22__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane6_strm1_data        ,
            output  wire                                        mgr22__std__lane6_strm1_data_valid  ,

            // manager 22, lane 7, stream 0      
            input   wire                                        std__mgr22__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane7_strm0_data        ,
            output  wire                                        mgr22__std__lane7_strm0_data_valid  ,

            // manager 22, lane 7, stream 1      
            input   wire                                        std__mgr22__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane7_strm1_data        ,
            output  wire                                        mgr22__std__lane7_strm1_data_valid  ,

            // manager 22, lane 8, stream 0      
            input   wire                                        std__mgr22__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane8_strm0_data        ,
            output  wire                                        mgr22__std__lane8_strm0_data_valid  ,

            // manager 22, lane 8, stream 1      
            input   wire                                        std__mgr22__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane8_strm1_data        ,
            output  wire                                        mgr22__std__lane8_strm1_data_valid  ,

            // manager 22, lane 9, stream 0      
            input   wire                                        std__mgr22__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane9_strm0_data        ,
            output  wire                                        mgr22__std__lane9_strm0_data_valid  ,

            // manager 22, lane 9, stream 1      
            input   wire                                        std__mgr22__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane9_strm1_data        ,
            output  wire                                        mgr22__std__lane9_strm1_data_valid  ,

            // manager 22, lane 10, stream 0      
            input   wire                                        std__mgr22__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane10_strm0_data        ,
            output  wire                                        mgr22__std__lane10_strm0_data_valid  ,

            // manager 22, lane 10, stream 1      
            input   wire                                        std__mgr22__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane10_strm1_data        ,
            output  wire                                        mgr22__std__lane10_strm1_data_valid  ,

            // manager 22, lane 11, stream 0      
            input   wire                                        std__mgr22__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane11_strm0_data        ,
            output  wire                                        mgr22__std__lane11_strm0_data_valid  ,

            // manager 22, lane 11, stream 1      
            input   wire                                        std__mgr22__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane11_strm1_data        ,
            output  wire                                        mgr22__std__lane11_strm1_data_valid  ,

            // manager 22, lane 12, stream 0      
            input   wire                                        std__mgr22__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane12_strm0_data        ,
            output  wire                                        mgr22__std__lane12_strm0_data_valid  ,

            // manager 22, lane 12, stream 1      
            input   wire                                        std__mgr22__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane12_strm1_data        ,
            output  wire                                        mgr22__std__lane12_strm1_data_valid  ,

            // manager 22, lane 13, stream 0      
            input   wire                                        std__mgr22__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane13_strm0_data        ,
            output  wire                                        mgr22__std__lane13_strm0_data_valid  ,

            // manager 22, lane 13, stream 1      
            input   wire                                        std__mgr22__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane13_strm1_data        ,
            output  wire                                        mgr22__std__lane13_strm1_data_valid  ,

            // manager 22, lane 14, stream 0      
            input   wire                                        std__mgr22__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane14_strm0_data        ,
            output  wire                                        mgr22__std__lane14_strm0_data_valid  ,

            // manager 22, lane 14, stream 1      
            input   wire                                        std__mgr22__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane14_strm1_data        ,
            output  wire                                        mgr22__std__lane14_strm1_data_valid  ,

            // manager 22, lane 15, stream 0      
            input   wire                                        std__mgr22__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane15_strm0_data        ,
            output  wire                                        mgr22__std__lane15_strm0_data_valid  ,

            // manager 22, lane 15, stream 1      
            input   wire                                        std__mgr22__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane15_strm1_data        ,
            output  wire                                        mgr22__std__lane15_strm1_data_valid  ,

            // manager 22, lane 16, stream 0      
            input   wire                                        std__mgr22__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane16_strm0_data        ,
            output  wire                                        mgr22__std__lane16_strm0_data_valid  ,

            // manager 22, lane 16, stream 1      
            input   wire                                        std__mgr22__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane16_strm1_data        ,
            output  wire                                        mgr22__std__lane16_strm1_data_valid  ,

            // manager 22, lane 17, stream 0      
            input   wire                                        std__mgr22__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane17_strm0_data        ,
            output  wire                                        mgr22__std__lane17_strm0_data_valid  ,

            // manager 22, lane 17, stream 1      
            input   wire                                        std__mgr22__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane17_strm1_data        ,
            output  wire                                        mgr22__std__lane17_strm1_data_valid  ,

            // manager 22, lane 18, stream 0      
            input   wire                                        std__mgr22__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane18_strm0_data        ,
            output  wire                                        mgr22__std__lane18_strm0_data_valid  ,

            // manager 22, lane 18, stream 1      
            input   wire                                        std__mgr22__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane18_strm1_data        ,
            output  wire                                        mgr22__std__lane18_strm1_data_valid  ,

            // manager 22, lane 19, stream 0      
            input   wire                                        std__mgr22__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane19_strm0_data        ,
            output  wire                                        mgr22__std__lane19_strm0_data_valid  ,

            // manager 22, lane 19, stream 1      
            input   wire                                        std__mgr22__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane19_strm1_data        ,
            output  wire                                        mgr22__std__lane19_strm1_data_valid  ,

            // manager 22, lane 20, stream 0      
            input   wire                                        std__mgr22__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane20_strm0_data        ,
            output  wire                                        mgr22__std__lane20_strm0_data_valid  ,

            // manager 22, lane 20, stream 1      
            input   wire                                        std__mgr22__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane20_strm1_data        ,
            output  wire                                        mgr22__std__lane20_strm1_data_valid  ,

            // manager 22, lane 21, stream 0      
            input   wire                                        std__mgr22__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane21_strm0_data        ,
            output  wire                                        mgr22__std__lane21_strm0_data_valid  ,

            // manager 22, lane 21, stream 1      
            input   wire                                        std__mgr22__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane21_strm1_data        ,
            output  wire                                        mgr22__std__lane21_strm1_data_valid  ,

            // manager 22, lane 22, stream 0      
            input   wire                                        std__mgr22__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane22_strm0_data        ,
            output  wire                                        mgr22__std__lane22_strm0_data_valid  ,

            // manager 22, lane 22, stream 1      
            input   wire                                        std__mgr22__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane22_strm1_data        ,
            output  wire                                        mgr22__std__lane22_strm1_data_valid  ,

            // manager 22, lane 23, stream 0      
            input   wire                                        std__mgr22__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane23_strm0_data        ,
            output  wire                                        mgr22__std__lane23_strm0_data_valid  ,

            // manager 22, lane 23, stream 1      
            input   wire                                        std__mgr22__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane23_strm1_data        ,
            output  wire                                        mgr22__std__lane23_strm1_data_valid  ,

            // manager 22, lane 24, stream 0      
            input   wire                                        std__mgr22__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane24_strm0_data        ,
            output  wire                                        mgr22__std__lane24_strm0_data_valid  ,

            // manager 22, lane 24, stream 1      
            input   wire                                        std__mgr22__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane24_strm1_data        ,
            output  wire                                        mgr22__std__lane24_strm1_data_valid  ,

            // manager 22, lane 25, stream 0      
            input   wire                                        std__mgr22__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane25_strm0_data        ,
            output  wire                                        mgr22__std__lane25_strm0_data_valid  ,

            // manager 22, lane 25, stream 1      
            input   wire                                        std__mgr22__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane25_strm1_data        ,
            output  wire                                        mgr22__std__lane25_strm1_data_valid  ,

            // manager 22, lane 26, stream 0      
            input   wire                                        std__mgr22__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane26_strm0_data        ,
            output  wire                                        mgr22__std__lane26_strm0_data_valid  ,

            // manager 22, lane 26, stream 1      
            input   wire                                        std__mgr22__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane26_strm1_data        ,
            output  wire                                        mgr22__std__lane26_strm1_data_valid  ,

            // manager 22, lane 27, stream 0      
            input   wire                                        std__mgr22__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane27_strm0_data        ,
            output  wire                                        mgr22__std__lane27_strm0_data_valid  ,

            // manager 22, lane 27, stream 1      
            input   wire                                        std__mgr22__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane27_strm1_data        ,
            output  wire                                        mgr22__std__lane27_strm1_data_valid  ,

            // manager 22, lane 28, stream 0      
            input   wire                                        std__mgr22__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane28_strm0_data        ,
            output  wire                                        mgr22__std__lane28_strm0_data_valid  ,

            // manager 22, lane 28, stream 1      
            input   wire                                        std__mgr22__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane28_strm1_data        ,
            output  wire                                        mgr22__std__lane28_strm1_data_valid  ,

            // manager 22, lane 29, stream 0      
            input   wire                                        std__mgr22__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane29_strm0_data        ,
            output  wire                                        mgr22__std__lane29_strm0_data_valid  ,

            // manager 22, lane 29, stream 1      
            input   wire                                        std__mgr22__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane29_strm1_data        ,
            output  wire                                        mgr22__std__lane29_strm1_data_valid  ,

            // manager 22, lane 30, stream 0      
            input   wire                                        std__mgr22__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane30_strm0_data        ,
            output  wire                                        mgr22__std__lane30_strm0_data_valid  ,

            // manager 22, lane 30, stream 1      
            input   wire                                        std__mgr22__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane30_strm1_data        ,
            output  wire                                        mgr22__std__lane30_strm1_data_valid  ,

            // manager 22, lane 31, stream 0      
            input   wire                                        std__mgr22__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane31_strm0_data        ,
            output  wire                                        mgr22__std__lane31_strm0_data_valid  ,

            // manager 22, lane 31, stream 1      
            input   wire                                        std__mgr22__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr22__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr22__std__lane31_strm1_data        ,
            output  wire                                        mgr22__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 23, lane 0, stream 0      
            input   wire                                        std__mgr23__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane0_strm0_data        ,
            output  wire                                        mgr23__std__lane0_strm0_data_valid  ,

            // manager 23, lane 0, stream 1      
            input   wire                                        std__mgr23__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane0_strm1_data        ,
            output  wire                                        mgr23__std__lane0_strm1_data_valid  ,

            // manager 23, lane 1, stream 0      
            input   wire                                        std__mgr23__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane1_strm0_data        ,
            output  wire                                        mgr23__std__lane1_strm0_data_valid  ,

            // manager 23, lane 1, stream 1      
            input   wire                                        std__mgr23__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane1_strm1_data        ,
            output  wire                                        mgr23__std__lane1_strm1_data_valid  ,

            // manager 23, lane 2, stream 0      
            input   wire                                        std__mgr23__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane2_strm0_data        ,
            output  wire                                        mgr23__std__lane2_strm0_data_valid  ,

            // manager 23, lane 2, stream 1      
            input   wire                                        std__mgr23__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane2_strm1_data        ,
            output  wire                                        mgr23__std__lane2_strm1_data_valid  ,

            // manager 23, lane 3, stream 0      
            input   wire                                        std__mgr23__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane3_strm0_data        ,
            output  wire                                        mgr23__std__lane3_strm0_data_valid  ,

            // manager 23, lane 3, stream 1      
            input   wire                                        std__mgr23__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane3_strm1_data        ,
            output  wire                                        mgr23__std__lane3_strm1_data_valid  ,

            // manager 23, lane 4, stream 0      
            input   wire                                        std__mgr23__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane4_strm0_data        ,
            output  wire                                        mgr23__std__lane4_strm0_data_valid  ,

            // manager 23, lane 4, stream 1      
            input   wire                                        std__mgr23__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane4_strm1_data        ,
            output  wire                                        mgr23__std__lane4_strm1_data_valid  ,

            // manager 23, lane 5, stream 0      
            input   wire                                        std__mgr23__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane5_strm0_data        ,
            output  wire                                        mgr23__std__lane5_strm0_data_valid  ,

            // manager 23, lane 5, stream 1      
            input   wire                                        std__mgr23__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane5_strm1_data        ,
            output  wire                                        mgr23__std__lane5_strm1_data_valid  ,

            // manager 23, lane 6, stream 0      
            input   wire                                        std__mgr23__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane6_strm0_data        ,
            output  wire                                        mgr23__std__lane6_strm0_data_valid  ,

            // manager 23, lane 6, stream 1      
            input   wire                                        std__mgr23__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane6_strm1_data        ,
            output  wire                                        mgr23__std__lane6_strm1_data_valid  ,

            // manager 23, lane 7, stream 0      
            input   wire                                        std__mgr23__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane7_strm0_data        ,
            output  wire                                        mgr23__std__lane7_strm0_data_valid  ,

            // manager 23, lane 7, stream 1      
            input   wire                                        std__mgr23__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane7_strm1_data        ,
            output  wire                                        mgr23__std__lane7_strm1_data_valid  ,

            // manager 23, lane 8, stream 0      
            input   wire                                        std__mgr23__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane8_strm0_data        ,
            output  wire                                        mgr23__std__lane8_strm0_data_valid  ,

            // manager 23, lane 8, stream 1      
            input   wire                                        std__mgr23__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane8_strm1_data        ,
            output  wire                                        mgr23__std__lane8_strm1_data_valid  ,

            // manager 23, lane 9, stream 0      
            input   wire                                        std__mgr23__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane9_strm0_data        ,
            output  wire                                        mgr23__std__lane9_strm0_data_valid  ,

            // manager 23, lane 9, stream 1      
            input   wire                                        std__mgr23__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane9_strm1_data        ,
            output  wire                                        mgr23__std__lane9_strm1_data_valid  ,

            // manager 23, lane 10, stream 0      
            input   wire                                        std__mgr23__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane10_strm0_data        ,
            output  wire                                        mgr23__std__lane10_strm0_data_valid  ,

            // manager 23, lane 10, stream 1      
            input   wire                                        std__mgr23__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane10_strm1_data        ,
            output  wire                                        mgr23__std__lane10_strm1_data_valid  ,

            // manager 23, lane 11, stream 0      
            input   wire                                        std__mgr23__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane11_strm0_data        ,
            output  wire                                        mgr23__std__lane11_strm0_data_valid  ,

            // manager 23, lane 11, stream 1      
            input   wire                                        std__mgr23__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane11_strm1_data        ,
            output  wire                                        mgr23__std__lane11_strm1_data_valid  ,

            // manager 23, lane 12, stream 0      
            input   wire                                        std__mgr23__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane12_strm0_data        ,
            output  wire                                        mgr23__std__lane12_strm0_data_valid  ,

            // manager 23, lane 12, stream 1      
            input   wire                                        std__mgr23__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane12_strm1_data        ,
            output  wire                                        mgr23__std__lane12_strm1_data_valid  ,

            // manager 23, lane 13, stream 0      
            input   wire                                        std__mgr23__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane13_strm0_data        ,
            output  wire                                        mgr23__std__lane13_strm0_data_valid  ,

            // manager 23, lane 13, stream 1      
            input   wire                                        std__mgr23__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane13_strm1_data        ,
            output  wire                                        mgr23__std__lane13_strm1_data_valid  ,

            // manager 23, lane 14, stream 0      
            input   wire                                        std__mgr23__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane14_strm0_data        ,
            output  wire                                        mgr23__std__lane14_strm0_data_valid  ,

            // manager 23, lane 14, stream 1      
            input   wire                                        std__mgr23__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane14_strm1_data        ,
            output  wire                                        mgr23__std__lane14_strm1_data_valid  ,

            // manager 23, lane 15, stream 0      
            input   wire                                        std__mgr23__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane15_strm0_data        ,
            output  wire                                        mgr23__std__lane15_strm0_data_valid  ,

            // manager 23, lane 15, stream 1      
            input   wire                                        std__mgr23__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane15_strm1_data        ,
            output  wire                                        mgr23__std__lane15_strm1_data_valid  ,

            // manager 23, lane 16, stream 0      
            input   wire                                        std__mgr23__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane16_strm0_data        ,
            output  wire                                        mgr23__std__lane16_strm0_data_valid  ,

            // manager 23, lane 16, stream 1      
            input   wire                                        std__mgr23__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane16_strm1_data        ,
            output  wire                                        mgr23__std__lane16_strm1_data_valid  ,

            // manager 23, lane 17, stream 0      
            input   wire                                        std__mgr23__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane17_strm0_data        ,
            output  wire                                        mgr23__std__lane17_strm0_data_valid  ,

            // manager 23, lane 17, stream 1      
            input   wire                                        std__mgr23__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane17_strm1_data        ,
            output  wire                                        mgr23__std__lane17_strm1_data_valid  ,

            // manager 23, lane 18, stream 0      
            input   wire                                        std__mgr23__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane18_strm0_data        ,
            output  wire                                        mgr23__std__lane18_strm0_data_valid  ,

            // manager 23, lane 18, stream 1      
            input   wire                                        std__mgr23__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane18_strm1_data        ,
            output  wire                                        mgr23__std__lane18_strm1_data_valid  ,

            // manager 23, lane 19, stream 0      
            input   wire                                        std__mgr23__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane19_strm0_data        ,
            output  wire                                        mgr23__std__lane19_strm0_data_valid  ,

            // manager 23, lane 19, stream 1      
            input   wire                                        std__mgr23__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane19_strm1_data        ,
            output  wire                                        mgr23__std__lane19_strm1_data_valid  ,

            // manager 23, lane 20, stream 0      
            input   wire                                        std__mgr23__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane20_strm0_data        ,
            output  wire                                        mgr23__std__lane20_strm0_data_valid  ,

            // manager 23, lane 20, stream 1      
            input   wire                                        std__mgr23__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane20_strm1_data        ,
            output  wire                                        mgr23__std__lane20_strm1_data_valid  ,

            // manager 23, lane 21, stream 0      
            input   wire                                        std__mgr23__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane21_strm0_data        ,
            output  wire                                        mgr23__std__lane21_strm0_data_valid  ,

            // manager 23, lane 21, stream 1      
            input   wire                                        std__mgr23__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane21_strm1_data        ,
            output  wire                                        mgr23__std__lane21_strm1_data_valid  ,

            // manager 23, lane 22, stream 0      
            input   wire                                        std__mgr23__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane22_strm0_data        ,
            output  wire                                        mgr23__std__lane22_strm0_data_valid  ,

            // manager 23, lane 22, stream 1      
            input   wire                                        std__mgr23__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane22_strm1_data        ,
            output  wire                                        mgr23__std__lane22_strm1_data_valid  ,

            // manager 23, lane 23, stream 0      
            input   wire                                        std__mgr23__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane23_strm0_data        ,
            output  wire                                        mgr23__std__lane23_strm0_data_valid  ,

            // manager 23, lane 23, stream 1      
            input   wire                                        std__mgr23__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane23_strm1_data        ,
            output  wire                                        mgr23__std__lane23_strm1_data_valid  ,

            // manager 23, lane 24, stream 0      
            input   wire                                        std__mgr23__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane24_strm0_data        ,
            output  wire                                        mgr23__std__lane24_strm0_data_valid  ,

            // manager 23, lane 24, stream 1      
            input   wire                                        std__mgr23__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane24_strm1_data        ,
            output  wire                                        mgr23__std__lane24_strm1_data_valid  ,

            // manager 23, lane 25, stream 0      
            input   wire                                        std__mgr23__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane25_strm0_data        ,
            output  wire                                        mgr23__std__lane25_strm0_data_valid  ,

            // manager 23, lane 25, stream 1      
            input   wire                                        std__mgr23__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane25_strm1_data        ,
            output  wire                                        mgr23__std__lane25_strm1_data_valid  ,

            // manager 23, lane 26, stream 0      
            input   wire                                        std__mgr23__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane26_strm0_data        ,
            output  wire                                        mgr23__std__lane26_strm0_data_valid  ,

            // manager 23, lane 26, stream 1      
            input   wire                                        std__mgr23__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane26_strm1_data        ,
            output  wire                                        mgr23__std__lane26_strm1_data_valid  ,

            // manager 23, lane 27, stream 0      
            input   wire                                        std__mgr23__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane27_strm0_data        ,
            output  wire                                        mgr23__std__lane27_strm0_data_valid  ,

            // manager 23, lane 27, stream 1      
            input   wire                                        std__mgr23__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane27_strm1_data        ,
            output  wire                                        mgr23__std__lane27_strm1_data_valid  ,

            // manager 23, lane 28, stream 0      
            input   wire                                        std__mgr23__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane28_strm0_data        ,
            output  wire                                        mgr23__std__lane28_strm0_data_valid  ,

            // manager 23, lane 28, stream 1      
            input   wire                                        std__mgr23__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane28_strm1_data        ,
            output  wire                                        mgr23__std__lane28_strm1_data_valid  ,

            // manager 23, lane 29, stream 0      
            input   wire                                        std__mgr23__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane29_strm0_data        ,
            output  wire                                        mgr23__std__lane29_strm0_data_valid  ,

            // manager 23, lane 29, stream 1      
            input   wire                                        std__mgr23__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane29_strm1_data        ,
            output  wire                                        mgr23__std__lane29_strm1_data_valid  ,

            // manager 23, lane 30, stream 0      
            input   wire                                        std__mgr23__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane30_strm0_data        ,
            output  wire                                        mgr23__std__lane30_strm0_data_valid  ,

            // manager 23, lane 30, stream 1      
            input   wire                                        std__mgr23__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane30_strm1_data        ,
            output  wire                                        mgr23__std__lane30_strm1_data_valid  ,

            // manager 23, lane 31, stream 0      
            input   wire                                        std__mgr23__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane31_strm0_data        ,
            output  wire                                        mgr23__std__lane31_strm0_data_valid  ,

            // manager 23, lane 31, stream 1      
            input   wire                                        std__mgr23__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr23__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr23__std__lane31_strm1_data        ,
            output  wire                                        mgr23__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 24, lane 0, stream 0      
            input   wire                                        std__mgr24__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane0_strm0_data        ,
            output  wire                                        mgr24__std__lane0_strm0_data_valid  ,

            // manager 24, lane 0, stream 1      
            input   wire                                        std__mgr24__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane0_strm1_data        ,
            output  wire                                        mgr24__std__lane0_strm1_data_valid  ,

            // manager 24, lane 1, stream 0      
            input   wire                                        std__mgr24__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane1_strm0_data        ,
            output  wire                                        mgr24__std__lane1_strm0_data_valid  ,

            // manager 24, lane 1, stream 1      
            input   wire                                        std__mgr24__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane1_strm1_data        ,
            output  wire                                        mgr24__std__lane1_strm1_data_valid  ,

            // manager 24, lane 2, stream 0      
            input   wire                                        std__mgr24__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane2_strm0_data        ,
            output  wire                                        mgr24__std__lane2_strm0_data_valid  ,

            // manager 24, lane 2, stream 1      
            input   wire                                        std__mgr24__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane2_strm1_data        ,
            output  wire                                        mgr24__std__lane2_strm1_data_valid  ,

            // manager 24, lane 3, stream 0      
            input   wire                                        std__mgr24__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane3_strm0_data        ,
            output  wire                                        mgr24__std__lane3_strm0_data_valid  ,

            // manager 24, lane 3, stream 1      
            input   wire                                        std__mgr24__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane3_strm1_data        ,
            output  wire                                        mgr24__std__lane3_strm1_data_valid  ,

            // manager 24, lane 4, stream 0      
            input   wire                                        std__mgr24__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane4_strm0_data        ,
            output  wire                                        mgr24__std__lane4_strm0_data_valid  ,

            // manager 24, lane 4, stream 1      
            input   wire                                        std__mgr24__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane4_strm1_data        ,
            output  wire                                        mgr24__std__lane4_strm1_data_valid  ,

            // manager 24, lane 5, stream 0      
            input   wire                                        std__mgr24__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane5_strm0_data        ,
            output  wire                                        mgr24__std__lane5_strm0_data_valid  ,

            // manager 24, lane 5, stream 1      
            input   wire                                        std__mgr24__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane5_strm1_data        ,
            output  wire                                        mgr24__std__lane5_strm1_data_valid  ,

            // manager 24, lane 6, stream 0      
            input   wire                                        std__mgr24__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane6_strm0_data        ,
            output  wire                                        mgr24__std__lane6_strm0_data_valid  ,

            // manager 24, lane 6, stream 1      
            input   wire                                        std__mgr24__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane6_strm1_data        ,
            output  wire                                        mgr24__std__lane6_strm1_data_valid  ,

            // manager 24, lane 7, stream 0      
            input   wire                                        std__mgr24__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane7_strm0_data        ,
            output  wire                                        mgr24__std__lane7_strm0_data_valid  ,

            // manager 24, lane 7, stream 1      
            input   wire                                        std__mgr24__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane7_strm1_data        ,
            output  wire                                        mgr24__std__lane7_strm1_data_valid  ,

            // manager 24, lane 8, stream 0      
            input   wire                                        std__mgr24__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane8_strm0_data        ,
            output  wire                                        mgr24__std__lane8_strm0_data_valid  ,

            // manager 24, lane 8, stream 1      
            input   wire                                        std__mgr24__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane8_strm1_data        ,
            output  wire                                        mgr24__std__lane8_strm1_data_valid  ,

            // manager 24, lane 9, stream 0      
            input   wire                                        std__mgr24__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane9_strm0_data        ,
            output  wire                                        mgr24__std__lane9_strm0_data_valid  ,

            // manager 24, lane 9, stream 1      
            input   wire                                        std__mgr24__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane9_strm1_data        ,
            output  wire                                        mgr24__std__lane9_strm1_data_valid  ,

            // manager 24, lane 10, stream 0      
            input   wire                                        std__mgr24__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane10_strm0_data        ,
            output  wire                                        mgr24__std__lane10_strm0_data_valid  ,

            // manager 24, lane 10, stream 1      
            input   wire                                        std__mgr24__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane10_strm1_data        ,
            output  wire                                        mgr24__std__lane10_strm1_data_valid  ,

            // manager 24, lane 11, stream 0      
            input   wire                                        std__mgr24__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane11_strm0_data        ,
            output  wire                                        mgr24__std__lane11_strm0_data_valid  ,

            // manager 24, lane 11, stream 1      
            input   wire                                        std__mgr24__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane11_strm1_data        ,
            output  wire                                        mgr24__std__lane11_strm1_data_valid  ,

            // manager 24, lane 12, stream 0      
            input   wire                                        std__mgr24__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane12_strm0_data        ,
            output  wire                                        mgr24__std__lane12_strm0_data_valid  ,

            // manager 24, lane 12, stream 1      
            input   wire                                        std__mgr24__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane12_strm1_data        ,
            output  wire                                        mgr24__std__lane12_strm1_data_valid  ,

            // manager 24, lane 13, stream 0      
            input   wire                                        std__mgr24__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane13_strm0_data        ,
            output  wire                                        mgr24__std__lane13_strm0_data_valid  ,

            // manager 24, lane 13, stream 1      
            input   wire                                        std__mgr24__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane13_strm1_data        ,
            output  wire                                        mgr24__std__lane13_strm1_data_valid  ,

            // manager 24, lane 14, stream 0      
            input   wire                                        std__mgr24__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane14_strm0_data        ,
            output  wire                                        mgr24__std__lane14_strm0_data_valid  ,

            // manager 24, lane 14, stream 1      
            input   wire                                        std__mgr24__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane14_strm1_data        ,
            output  wire                                        mgr24__std__lane14_strm1_data_valid  ,

            // manager 24, lane 15, stream 0      
            input   wire                                        std__mgr24__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane15_strm0_data        ,
            output  wire                                        mgr24__std__lane15_strm0_data_valid  ,

            // manager 24, lane 15, stream 1      
            input   wire                                        std__mgr24__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane15_strm1_data        ,
            output  wire                                        mgr24__std__lane15_strm1_data_valid  ,

            // manager 24, lane 16, stream 0      
            input   wire                                        std__mgr24__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane16_strm0_data        ,
            output  wire                                        mgr24__std__lane16_strm0_data_valid  ,

            // manager 24, lane 16, stream 1      
            input   wire                                        std__mgr24__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane16_strm1_data        ,
            output  wire                                        mgr24__std__lane16_strm1_data_valid  ,

            // manager 24, lane 17, stream 0      
            input   wire                                        std__mgr24__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane17_strm0_data        ,
            output  wire                                        mgr24__std__lane17_strm0_data_valid  ,

            // manager 24, lane 17, stream 1      
            input   wire                                        std__mgr24__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane17_strm1_data        ,
            output  wire                                        mgr24__std__lane17_strm1_data_valid  ,

            // manager 24, lane 18, stream 0      
            input   wire                                        std__mgr24__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane18_strm0_data        ,
            output  wire                                        mgr24__std__lane18_strm0_data_valid  ,

            // manager 24, lane 18, stream 1      
            input   wire                                        std__mgr24__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane18_strm1_data        ,
            output  wire                                        mgr24__std__lane18_strm1_data_valid  ,

            // manager 24, lane 19, stream 0      
            input   wire                                        std__mgr24__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane19_strm0_data        ,
            output  wire                                        mgr24__std__lane19_strm0_data_valid  ,

            // manager 24, lane 19, stream 1      
            input   wire                                        std__mgr24__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane19_strm1_data        ,
            output  wire                                        mgr24__std__lane19_strm1_data_valid  ,

            // manager 24, lane 20, stream 0      
            input   wire                                        std__mgr24__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane20_strm0_data        ,
            output  wire                                        mgr24__std__lane20_strm0_data_valid  ,

            // manager 24, lane 20, stream 1      
            input   wire                                        std__mgr24__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane20_strm1_data        ,
            output  wire                                        mgr24__std__lane20_strm1_data_valid  ,

            // manager 24, lane 21, stream 0      
            input   wire                                        std__mgr24__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane21_strm0_data        ,
            output  wire                                        mgr24__std__lane21_strm0_data_valid  ,

            // manager 24, lane 21, stream 1      
            input   wire                                        std__mgr24__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane21_strm1_data        ,
            output  wire                                        mgr24__std__lane21_strm1_data_valid  ,

            // manager 24, lane 22, stream 0      
            input   wire                                        std__mgr24__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane22_strm0_data        ,
            output  wire                                        mgr24__std__lane22_strm0_data_valid  ,

            // manager 24, lane 22, stream 1      
            input   wire                                        std__mgr24__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane22_strm1_data        ,
            output  wire                                        mgr24__std__lane22_strm1_data_valid  ,

            // manager 24, lane 23, stream 0      
            input   wire                                        std__mgr24__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane23_strm0_data        ,
            output  wire                                        mgr24__std__lane23_strm0_data_valid  ,

            // manager 24, lane 23, stream 1      
            input   wire                                        std__mgr24__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane23_strm1_data        ,
            output  wire                                        mgr24__std__lane23_strm1_data_valid  ,

            // manager 24, lane 24, stream 0      
            input   wire                                        std__mgr24__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane24_strm0_data        ,
            output  wire                                        mgr24__std__lane24_strm0_data_valid  ,

            // manager 24, lane 24, stream 1      
            input   wire                                        std__mgr24__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane24_strm1_data        ,
            output  wire                                        mgr24__std__lane24_strm1_data_valid  ,

            // manager 24, lane 25, stream 0      
            input   wire                                        std__mgr24__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane25_strm0_data        ,
            output  wire                                        mgr24__std__lane25_strm0_data_valid  ,

            // manager 24, lane 25, stream 1      
            input   wire                                        std__mgr24__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane25_strm1_data        ,
            output  wire                                        mgr24__std__lane25_strm1_data_valid  ,

            // manager 24, lane 26, stream 0      
            input   wire                                        std__mgr24__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane26_strm0_data        ,
            output  wire                                        mgr24__std__lane26_strm0_data_valid  ,

            // manager 24, lane 26, stream 1      
            input   wire                                        std__mgr24__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane26_strm1_data        ,
            output  wire                                        mgr24__std__lane26_strm1_data_valid  ,

            // manager 24, lane 27, stream 0      
            input   wire                                        std__mgr24__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane27_strm0_data        ,
            output  wire                                        mgr24__std__lane27_strm0_data_valid  ,

            // manager 24, lane 27, stream 1      
            input   wire                                        std__mgr24__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane27_strm1_data        ,
            output  wire                                        mgr24__std__lane27_strm1_data_valid  ,

            // manager 24, lane 28, stream 0      
            input   wire                                        std__mgr24__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane28_strm0_data        ,
            output  wire                                        mgr24__std__lane28_strm0_data_valid  ,

            // manager 24, lane 28, stream 1      
            input   wire                                        std__mgr24__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane28_strm1_data        ,
            output  wire                                        mgr24__std__lane28_strm1_data_valid  ,

            // manager 24, lane 29, stream 0      
            input   wire                                        std__mgr24__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane29_strm0_data        ,
            output  wire                                        mgr24__std__lane29_strm0_data_valid  ,

            // manager 24, lane 29, stream 1      
            input   wire                                        std__mgr24__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane29_strm1_data        ,
            output  wire                                        mgr24__std__lane29_strm1_data_valid  ,

            // manager 24, lane 30, stream 0      
            input   wire                                        std__mgr24__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane30_strm0_data        ,
            output  wire                                        mgr24__std__lane30_strm0_data_valid  ,

            // manager 24, lane 30, stream 1      
            input   wire                                        std__mgr24__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane30_strm1_data        ,
            output  wire                                        mgr24__std__lane30_strm1_data_valid  ,

            // manager 24, lane 31, stream 0      
            input   wire                                        std__mgr24__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane31_strm0_data        ,
            output  wire                                        mgr24__std__lane31_strm0_data_valid  ,

            // manager 24, lane 31, stream 1      
            input   wire                                        std__mgr24__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr24__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr24__std__lane31_strm1_data        ,
            output  wire                                        mgr24__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 25, lane 0, stream 0      
            input   wire                                        std__mgr25__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane0_strm0_data        ,
            output  wire                                        mgr25__std__lane0_strm0_data_valid  ,

            // manager 25, lane 0, stream 1      
            input   wire                                        std__mgr25__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane0_strm1_data        ,
            output  wire                                        mgr25__std__lane0_strm1_data_valid  ,

            // manager 25, lane 1, stream 0      
            input   wire                                        std__mgr25__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane1_strm0_data        ,
            output  wire                                        mgr25__std__lane1_strm0_data_valid  ,

            // manager 25, lane 1, stream 1      
            input   wire                                        std__mgr25__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane1_strm1_data        ,
            output  wire                                        mgr25__std__lane1_strm1_data_valid  ,

            // manager 25, lane 2, stream 0      
            input   wire                                        std__mgr25__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane2_strm0_data        ,
            output  wire                                        mgr25__std__lane2_strm0_data_valid  ,

            // manager 25, lane 2, stream 1      
            input   wire                                        std__mgr25__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane2_strm1_data        ,
            output  wire                                        mgr25__std__lane2_strm1_data_valid  ,

            // manager 25, lane 3, stream 0      
            input   wire                                        std__mgr25__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane3_strm0_data        ,
            output  wire                                        mgr25__std__lane3_strm0_data_valid  ,

            // manager 25, lane 3, stream 1      
            input   wire                                        std__mgr25__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane3_strm1_data        ,
            output  wire                                        mgr25__std__lane3_strm1_data_valid  ,

            // manager 25, lane 4, stream 0      
            input   wire                                        std__mgr25__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane4_strm0_data        ,
            output  wire                                        mgr25__std__lane4_strm0_data_valid  ,

            // manager 25, lane 4, stream 1      
            input   wire                                        std__mgr25__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane4_strm1_data        ,
            output  wire                                        mgr25__std__lane4_strm1_data_valid  ,

            // manager 25, lane 5, stream 0      
            input   wire                                        std__mgr25__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane5_strm0_data        ,
            output  wire                                        mgr25__std__lane5_strm0_data_valid  ,

            // manager 25, lane 5, stream 1      
            input   wire                                        std__mgr25__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane5_strm1_data        ,
            output  wire                                        mgr25__std__lane5_strm1_data_valid  ,

            // manager 25, lane 6, stream 0      
            input   wire                                        std__mgr25__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane6_strm0_data        ,
            output  wire                                        mgr25__std__lane6_strm0_data_valid  ,

            // manager 25, lane 6, stream 1      
            input   wire                                        std__mgr25__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane6_strm1_data        ,
            output  wire                                        mgr25__std__lane6_strm1_data_valid  ,

            // manager 25, lane 7, stream 0      
            input   wire                                        std__mgr25__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane7_strm0_data        ,
            output  wire                                        mgr25__std__lane7_strm0_data_valid  ,

            // manager 25, lane 7, stream 1      
            input   wire                                        std__mgr25__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane7_strm1_data        ,
            output  wire                                        mgr25__std__lane7_strm1_data_valid  ,

            // manager 25, lane 8, stream 0      
            input   wire                                        std__mgr25__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane8_strm0_data        ,
            output  wire                                        mgr25__std__lane8_strm0_data_valid  ,

            // manager 25, lane 8, stream 1      
            input   wire                                        std__mgr25__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane8_strm1_data        ,
            output  wire                                        mgr25__std__lane8_strm1_data_valid  ,

            // manager 25, lane 9, stream 0      
            input   wire                                        std__mgr25__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane9_strm0_data        ,
            output  wire                                        mgr25__std__lane9_strm0_data_valid  ,

            // manager 25, lane 9, stream 1      
            input   wire                                        std__mgr25__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane9_strm1_data        ,
            output  wire                                        mgr25__std__lane9_strm1_data_valid  ,

            // manager 25, lane 10, stream 0      
            input   wire                                        std__mgr25__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane10_strm0_data        ,
            output  wire                                        mgr25__std__lane10_strm0_data_valid  ,

            // manager 25, lane 10, stream 1      
            input   wire                                        std__mgr25__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane10_strm1_data        ,
            output  wire                                        mgr25__std__lane10_strm1_data_valid  ,

            // manager 25, lane 11, stream 0      
            input   wire                                        std__mgr25__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane11_strm0_data        ,
            output  wire                                        mgr25__std__lane11_strm0_data_valid  ,

            // manager 25, lane 11, stream 1      
            input   wire                                        std__mgr25__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane11_strm1_data        ,
            output  wire                                        mgr25__std__lane11_strm1_data_valid  ,

            // manager 25, lane 12, stream 0      
            input   wire                                        std__mgr25__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane12_strm0_data        ,
            output  wire                                        mgr25__std__lane12_strm0_data_valid  ,

            // manager 25, lane 12, stream 1      
            input   wire                                        std__mgr25__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane12_strm1_data        ,
            output  wire                                        mgr25__std__lane12_strm1_data_valid  ,

            // manager 25, lane 13, stream 0      
            input   wire                                        std__mgr25__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane13_strm0_data        ,
            output  wire                                        mgr25__std__lane13_strm0_data_valid  ,

            // manager 25, lane 13, stream 1      
            input   wire                                        std__mgr25__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane13_strm1_data        ,
            output  wire                                        mgr25__std__lane13_strm1_data_valid  ,

            // manager 25, lane 14, stream 0      
            input   wire                                        std__mgr25__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane14_strm0_data        ,
            output  wire                                        mgr25__std__lane14_strm0_data_valid  ,

            // manager 25, lane 14, stream 1      
            input   wire                                        std__mgr25__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane14_strm1_data        ,
            output  wire                                        mgr25__std__lane14_strm1_data_valid  ,

            // manager 25, lane 15, stream 0      
            input   wire                                        std__mgr25__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane15_strm0_data        ,
            output  wire                                        mgr25__std__lane15_strm0_data_valid  ,

            // manager 25, lane 15, stream 1      
            input   wire                                        std__mgr25__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane15_strm1_data        ,
            output  wire                                        mgr25__std__lane15_strm1_data_valid  ,

            // manager 25, lane 16, stream 0      
            input   wire                                        std__mgr25__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane16_strm0_data        ,
            output  wire                                        mgr25__std__lane16_strm0_data_valid  ,

            // manager 25, lane 16, stream 1      
            input   wire                                        std__mgr25__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane16_strm1_data        ,
            output  wire                                        mgr25__std__lane16_strm1_data_valid  ,

            // manager 25, lane 17, stream 0      
            input   wire                                        std__mgr25__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane17_strm0_data        ,
            output  wire                                        mgr25__std__lane17_strm0_data_valid  ,

            // manager 25, lane 17, stream 1      
            input   wire                                        std__mgr25__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane17_strm1_data        ,
            output  wire                                        mgr25__std__lane17_strm1_data_valid  ,

            // manager 25, lane 18, stream 0      
            input   wire                                        std__mgr25__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane18_strm0_data        ,
            output  wire                                        mgr25__std__lane18_strm0_data_valid  ,

            // manager 25, lane 18, stream 1      
            input   wire                                        std__mgr25__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane18_strm1_data        ,
            output  wire                                        mgr25__std__lane18_strm1_data_valid  ,

            // manager 25, lane 19, stream 0      
            input   wire                                        std__mgr25__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane19_strm0_data        ,
            output  wire                                        mgr25__std__lane19_strm0_data_valid  ,

            // manager 25, lane 19, stream 1      
            input   wire                                        std__mgr25__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane19_strm1_data        ,
            output  wire                                        mgr25__std__lane19_strm1_data_valid  ,

            // manager 25, lane 20, stream 0      
            input   wire                                        std__mgr25__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane20_strm0_data        ,
            output  wire                                        mgr25__std__lane20_strm0_data_valid  ,

            // manager 25, lane 20, stream 1      
            input   wire                                        std__mgr25__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane20_strm1_data        ,
            output  wire                                        mgr25__std__lane20_strm1_data_valid  ,

            // manager 25, lane 21, stream 0      
            input   wire                                        std__mgr25__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane21_strm0_data        ,
            output  wire                                        mgr25__std__lane21_strm0_data_valid  ,

            // manager 25, lane 21, stream 1      
            input   wire                                        std__mgr25__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane21_strm1_data        ,
            output  wire                                        mgr25__std__lane21_strm1_data_valid  ,

            // manager 25, lane 22, stream 0      
            input   wire                                        std__mgr25__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane22_strm0_data        ,
            output  wire                                        mgr25__std__lane22_strm0_data_valid  ,

            // manager 25, lane 22, stream 1      
            input   wire                                        std__mgr25__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane22_strm1_data        ,
            output  wire                                        mgr25__std__lane22_strm1_data_valid  ,

            // manager 25, lane 23, stream 0      
            input   wire                                        std__mgr25__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane23_strm0_data        ,
            output  wire                                        mgr25__std__lane23_strm0_data_valid  ,

            // manager 25, lane 23, stream 1      
            input   wire                                        std__mgr25__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane23_strm1_data        ,
            output  wire                                        mgr25__std__lane23_strm1_data_valid  ,

            // manager 25, lane 24, stream 0      
            input   wire                                        std__mgr25__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane24_strm0_data        ,
            output  wire                                        mgr25__std__lane24_strm0_data_valid  ,

            // manager 25, lane 24, stream 1      
            input   wire                                        std__mgr25__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane24_strm1_data        ,
            output  wire                                        mgr25__std__lane24_strm1_data_valid  ,

            // manager 25, lane 25, stream 0      
            input   wire                                        std__mgr25__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane25_strm0_data        ,
            output  wire                                        mgr25__std__lane25_strm0_data_valid  ,

            // manager 25, lane 25, stream 1      
            input   wire                                        std__mgr25__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane25_strm1_data        ,
            output  wire                                        mgr25__std__lane25_strm1_data_valid  ,

            // manager 25, lane 26, stream 0      
            input   wire                                        std__mgr25__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane26_strm0_data        ,
            output  wire                                        mgr25__std__lane26_strm0_data_valid  ,

            // manager 25, lane 26, stream 1      
            input   wire                                        std__mgr25__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane26_strm1_data        ,
            output  wire                                        mgr25__std__lane26_strm1_data_valid  ,

            // manager 25, lane 27, stream 0      
            input   wire                                        std__mgr25__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane27_strm0_data        ,
            output  wire                                        mgr25__std__lane27_strm0_data_valid  ,

            // manager 25, lane 27, stream 1      
            input   wire                                        std__mgr25__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane27_strm1_data        ,
            output  wire                                        mgr25__std__lane27_strm1_data_valid  ,

            // manager 25, lane 28, stream 0      
            input   wire                                        std__mgr25__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane28_strm0_data        ,
            output  wire                                        mgr25__std__lane28_strm0_data_valid  ,

            // manager 25, lane 28, stream 1      
            input   wire                                        std__mgr25__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane28_strm1_data        ,
            output  wire                                        mgr25__std__lane28_strm1_data_valid  ,

            // manager 25, lane 29, stream 0      
            input   wire                                        std__mgr25__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane29_strm0_data        ,
            output  wire                                        mgr25__std__lane29_strm0_data_valid  ,

            // manager 25, lane 29, stream 1      
            input   wire                                        std__mgr25__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane29_strm1_data        ,
            output  wire                                        mgr25__std__lane29_strm1_data_valid  ,

            // manager 25, lane 30, stream 0      
            input   wire                                        std__mgr25__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane30_strm0_data        ,
            output  wire                                        mgr25__std__lane30_strm0_data_valid  ,

            // manager 25, lane 30, stream 1      
            input   wire                                        std__mgr25__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane30_strm1_data        ,
            output  wire                                        mgr25__std__lane30_strm1_data_valid  ,

            // manager 25, lane 31, stream 0      
            input   wire                                        std__mgr25__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane31_strm0_data        ,
            output  wire                                        mgr25__std__lane31_strm0_data_valid  ,

            // manager 25, lane 31, stream 1      
            input   wire                                        std__mgr25__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr25__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr25__std__lane31_strm1_data        ,
            output  wire                                        mgr25__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 26, lane 0, stream 0      
            input   wire                                        std__mgr26__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane0_strm0_data        ,
            output  wire                                        mgr26__std__lane0_strm0_data_valid  ,

            // manager 26, lane 0, stream 1      
            input   wire                                        std__mgr26__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane0_strm1_data        ,
            output  wire                                        mgr26__std__lane0_strm1_data_valid  ,

            // manager 26, lane 1, stream 0      
            input   wire                                        std__mgr26__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane1_strm0_data        ,
            output  wire                                        mgr26__std__lane1_strm0_data_valid  ,

            // manager 26, lane 1, stream 1      
            input   wire                                        std__mgr26__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane1_strm1_data        ,
            output  wire                                        mgr26__std__lane1_strm1_data_valid  ,

            // manager 26, lane 2, stream 0      
            input   wire                                        std__mgr26__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane2_strm0_data        ,
            output  wire                                        mgr26__std__lane2_strm0_data_valid  ,

            // manager 26, lane 2, stream 1      
            input   wire                                        std__mgr26__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane2_strm1_data        ,
            output  wire                                        mgr26__std__lane2_strm1_data_valid  ,

            // manager 26, lane 3, stream 0      
            input   wire                                        std__mgr26__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane3_strm0_data        ,
            output  wire                                        mgr26__std__lane3_strm0_data_valid  ,

            // manager 26, lane 3, stream 1      
            input   wire                                        std__mgr26__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane3_strm1_data        ,
            output  wire                                        mgr26__std__lane3_strm1_data_valid  ,

            // manager 26, lane 4, stream 0      
            input   wire                                        std__mgr26__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane4_strm0_data        ,
            output  wire                                        mgr26__std__lane4_strm0_data_valid  ,

            // manager 26, lane 4, stream 1      
            input   wire                                        std__mgr26__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane4_strm1_data        ,
            output  wire                                        mgr26__std__lane4_strm1_data_valid  ,

            // manager 26, lane 5, stream 0      
            input   wire                                        std__mgr26__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane5_strm0_data        ,
            output  wire                                        mgr26__std__lane5_strm0_data_valid  ,

            // manager 26, lane 5, stream 1      
            input   wire                                        std__mgr26__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane5_strm1_data        ,
            output  wire                                        mgr26__std__lane5_strm1_data_valid  ,

            // manager 26, lane 6, stream 0      
            input   wire                                        std__mgr26__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane6_strm0_data        ,
            output  wire                                        mgr26__std__lane6_strm0_data_valid  ,

            // manager 26, lane 6, stream 1      
            input   wire                                        std__mgr26__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane6_strm1_data        ,
            output  wire                                        mgr26__std__lane6_strm1_data_valid  ,

            // manager 26, lane 7, stream 0      
            input   wire                                        std__mgr26__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane7_strm0_data        ,
            output  wire                                        mgr26__std__lane7_strm0_data_valid  ,

            // manager 26, lane 7, stream 1      
            input   wire                                        std__mgr26__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane7_strm1_data        ,
            output  wire                                        mgr26__std__lane7_strm1_data_valid  ,

            // manager 26, lane 8, stream 0      
            input   wire                                        std__mgr26__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane8_strm0_data        ,
            output  wire                                        mgr26__std__lane8_strm0_data_valid  ,

            // manager 26, lane 8, stream 1      
            input   wire                                        std__mgr26__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane8_strm1_data        ,
            output  wire                                        mgr26__std__lane8_strm1_data_valid  ,

            // manager 26, lane 9, stream 0      
            input   wire                                        std__mgr26__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane9_strm0_data        ,
            output  wire                                        mgr26__std__lane9_strm0_data_valid  ,

            // manager 26, lane 9, stream 1      
            input   wire                                        std__mgr26__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane9_strm1_data        ,
            output  wire                                        mgr26__std__lane9_strm1_data_valid  ,

            // manager 26, lane 10, stream 0      
            input   wire                                        std__mgr26__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane10_strm0_data        ,
            output  wire                                        mgr26__std__lane10_strm0_data_valid  ,

            // manager 26, lane 10, stream 1      
            input   wire                                        std__mgr26__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane10_strm1_data        ,
            output  wire                                        mgr26__std__lane10_strm1_data_valid  ,

            // manager 26, lane 11, stream 0      
            input   wire                                        std__mgr26__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane11_strm0_data        ,
            output  wire                                        mgr26__std__lane11_strm0_data_valid  ,

            // manager 26, lane 11, stream 1      
            input   wire                                        std__mgr26__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane11_strm1_data        ,
            output  wire                                        mgr26__std__lane11_strm1_data_valid  ,

            // manager 26, lane 12, stream 0      
            input   wire                                        std__mgr26__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane12_strm0_data        ,
            output  wire                                        mgr26__std__lane12_strm0_data_valid  ,

            // manager 26, lane 12, stream 1      
            input   wire                                        std__mgr26__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane12_strm1_data        ,
            output  wire                                        mgr26__std__lane12_strm1_data_valid  ,

            // manager 26, lane 13, stream 0      
            input   wire                                        std__mgr26__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane13_strm0_data        ,
            output  wire                                        mgr26__std__lane13_strm0_data_valid  ,

            // manager 26, lane 13, stream 1      
            input   wire                                        std__mgr26__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane13_strm1_data        ,
            output  wire                                        mgr26__std__lane13_strm1_data_valid  ,

            // manager 26, lane 14, stream 0      
            input   wire                                        std__mgr26__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane14_strm0_data        ,
            output  wire                                        mgr26__std__lane14_strm0_data_valid  ,

            // manager 26, lane 14, stream 1      
            input   wire                                        std__mgr26__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane14_strm1_data        ,
            output  wire                                        mgr26__std__lane14_strm1_data_valid  ,

            // manager 26, lane 15, stream 0      
            input   wire                                        std__mgr26__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane15_strm0_data        ,
            output  wire                                        mgr26__std__lane15_strm0_data_valid  ,

            // manager 26, lane 15, stream 1      
            input   wire                                        std__mgr26__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane15_strm1_data        ,
            output  wire                                        mgr26__std__lane15_strm1_data_valid  ,

            // manager 26, lane 16, stream 0      
            input   wire                                        std__mgr26__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane16_strm0_data        ,
            output  wire                                        mgr26__std__lane16_strm0_data_valid  ,

            // manager 26, lane 16, stream 1      
            input   wire                                        std__mgr26__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane16_strm1_data        ,
            output  wire                                        mgr26__std__lane16_strm1_data_valid  ,

            // manager 26, lane 17, stream 0      
            input   wire                                        std__mgr26__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane17_strm0_data        ,
            output  wire                                        mgr26__std__lane17_strm0_data_valid  ,

            // manager 26, lane 17, stream 1      
            input   wire                                        std__mgr26__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane17_strm1_data        ,
            output  wire                                        mgr26__std__lane17_strm1_data_valid  ,

            // manager 26, lane 18, stream 0      
            input   wire                                        std__mgr26__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane18_strm0_data        ,
            output  wire                                        mgr26__std__lane18_strm0_data_valid  ,

            // manager 26, lane 18, stream 1      
            input   wire                                        std__mgr26__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane18_strm1_data        ,
            output  wire                                        mgr26__std__lane18_strm1_data_valid  ,

            // manager 26, lane 19, stream 0      
            input   wire                                        std__mgr26__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane19_strm0_data        ,
            output  wire                                        mgr26__std__lane19_strm0_data_valid  ,

            // manager 26, lane 19, stream 1      
            input   wire                                        std__mgr26__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane19_strm1_data        ,
            output  wire                                        mgr26__std__lane19_strm1_data_valid  ,

            // manager 26, lane 20, stream 0      
            input   wire                                        std__mgr26__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane20_strm0_data        ,
            output  wire                                        mgr26__std__lane20_strm0_data_valid  ,

            // manager 26, lane 20, stream 1      
            input   wire                                        std__mgr26__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane20_strm1_data        ,
            output  wire                                        mgr26__std__lane20_strm1_data_valid  ,

            // manager 26, lane 21, stream 0      
            input   wire                                        std__mgr26__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane21_strm0_data        ,
            output  wire                                        mgr26__std__lane21_strm0_data_valid  ,

            // manager 26, lane 21, stream 1      
            input   wire                                        std__mgr26__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane21_strm1_data        ,
            output  wire                                        mgr26__std__lane21_strm1_data_valid  ,

            // manager 26, lane 22, stream 0      
            input   wire                                        std__mgr26__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane22_strm0_data        ,
            output  wire                                        mgr26__std__lane22_strm0_data_valid  ,

            // manager 26, lane 22, stream 1      
            input   wire                                        std__mgr26__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane22_strm1_data        ,
            output  wire                                        mgr26__std__lane22_strm1_data_valid  ,

            // manager 26, lane 23, stream 0      
            input   wire                                        std__mgr26__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane23_strm0_data        ,
            output  wire                                        mgr26__std__lane23_strm0_data_valid  ,

            // manager 26, lane 23, stream 1      
            input   wire                                        std__mgr26__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane23_strm1_data        ,
            output  wire                                        mgr26__std__lane23_strm1_data_valid  ,

            // manager 26, lane 24, stream 0      
            input   wire                                        std__mgr26__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane24_strm0_data        ,
            output  wire                                        mgr26__std__lane24_strm0_data_valid  ,

            // manager 26, lane 24, stream 1      
            input   wire                                        std__mgr26__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane24_strm1_data        ,
            output  wire                                        mgr26__std__lane24_strm1_data_valid  ,

            // manager 26, lane 25, stream 0      
            input   wire                                        std__mgr26__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane25_strm0_data        ,
            output  wire                                        mgr26__std__lane25_strm0_data_valid  ,

            // manager 26, lane 25, stream 1      
            input   wire                                        std__mgr26__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane25_strm1_data        ,
            output  wire                                        mgr26__std__lane25_strm1_data_valid  ,

            // manager 26, lane 26, stream 0      
            input   wire                                        std__mgr26__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane26_strm0_data        ,
            output  wire                                        mgr26__std__lane26_strm0_data_valid  ,

            // manager 26, lane 26, stream 1      
            input   wire                                        std__mgr26__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane26_strm1_data        ,
            output  wire                                        mgr26__std__lane26_strm1_data_valid  ,

            // manager 26, lane 27, stream 0      
            input   wire                                        std__mgr26__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane27_strm0_data        ,
            output  wire                                        mgr26__std__lane27_strm0_data_valid  ,

            // manager 26, lane 27, stream 1      
            input   wire                                        std__mgr26__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane27_strm1_data        ,
            output  wire                                        mgr26__std__lane27_strm1_data_valid  ,

            // manager 26, lane 28, stream 0      
            input   wire                                        std__mgr26__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane28_strm0_data        ,
            output  wire                                        mgr26__std__lane28_strm0_data_valid  ,

            // manager 26, lane 28, stream 1      
            input   wire                                        std__mgr26__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane28_strm1_data        ,
            output  wire                                        mgr26__std__lane28_strm1_data_valid  ,

            // manager 26, lane 29, stream 0      
            input   wire                                        std__mgr26__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane29_strm0_data        ,
            output  wire                                        mgr26__std__lane29_strm0_data_valid  ,

            // manager 26, lane 29, stream 1      
            input   wire                                        std__mgr26__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane29_strm1_data        ,
            output  wire                                        mgr26__std__lane29_strm1_data_valid  ,

            // manager 26, lane 30, stream 0      
            input   wire                                        std__mgr26__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane30_strm0_data        ,
            output  wire                                        mgr26__std__lane30_strm0_data_valid  ,

            // manager 26, lane 30, stream 1      
            input   wire                                        std__mgr26__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane30_strm1_data        ,
            output  wire                                        mgr26__std__lane30_strm1_data_valid  ,

            // manager 26, lane 31, stream 0      
            input   wire                                        std__mgr26__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane31_strm0_data        ,
            output  wire                                        mgr26__std__lane31_strm0_data_valid  ,

            // manager 26, lane 31, stream 1      
            input   wire                                        std__mgr26__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr26__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr26__std__lane31_strm1_data        ,
            output  wire                                        mgr26__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 27, lane 0, stream 0      
            input   wire                                        std__mgr27__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane0_strm0_data        ,
            output  wire                                        mgr27__std__lane0_strm0_data_valid  ,

            // manager 27, lane 0, stream 1      
            input   wire                                        std__mgr27__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane0_strm1_data        ,
            output  wire                                        mgr27__std__lane0_strm1_data_valid  ,

            // manager 27, lane 1, stream 0      
            input   wire                                        std__mgr27__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane1_strm0_data        ,
            output  wire                                        mgr27__std__lane1_strm0_data_valid  ,

            // manager 27, lane 1, stream 1      
            input   wire                                        std__mgr27__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane1_strm1_data        ,
            output  wire                                        mgr27__std__lane1_strm1_data_valid  ,

            // manager 27, lane 2, stream 0      
            input   wire                                        std__mgr27__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane2_strm0_data        ,
            output  wire                                        mgr27__std__lane2_strm0_data_valid  ,

            // manager 27, lane 2, stream 1      
            input   wire                                        std__mgr27__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane2_strm1_data        ,
            output  wire                                        mgr27__std__lane2_strm1_data_valid  ,

            // manager 27, lane 3, stream 0      
            input   wire                                        std__mgr27__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane3_strm0_data        ,
            output  wire                                        mgr27__std__lane3_strm0_data_valid  ,

            // manager 27, lane 3, stream 1      
            input   wire                                        std__mgr27__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane3_strm1_data        ,
            output  wire                                        mgr27__std__lane3_strm1_data_valid  ,

            // manager 27, lane 4, stream 0      
            input   wire                                        std__mgr27__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane4_strm0_data        ,
            output  wire                                        mgr27__std__lane4_strm0_data_valid  ,

            // manager 27, lane 4, stream 1      
            input   wire                                        std__mgr27__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane4_strm1_data        ,
            output  wire                                        mgr27__std__lane4_strm1_data_valid  ,

            // manager 27, lane 5, stream 0      
            input   wire                                        std__mgr27__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane5_strm0_data        ,
            output  wire                                        mgr27__std__lane5_strm0_data_valid  ,

            // manager 27, lane 5, stream 1      
            input   wire                                        std__mgr27__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane5_strm1_data        ,
            output  wire                                        mgr27__std__lane5_strm1_data_valid  ,

            // manager 27, lane 6, stream 0      
            input   wire                                        std__mgr27__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane6_strm0_data        ,
            output  wire                                        mgr27__std__lane6_strm0_data_valid  ,

            // manager 27, lane 6, stream 1      
            input   wire                                        std__mgr27__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane6_strm1_data        ,
            output  wire                                        mgr27__std__lane6_strm1_data_valid  ,

            // manager 27, lane 7, stream 0      
            input   wire                                        std__mgr27__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane7_strm0_data        ,
            output  wire                                        mgr27__std__lane7_strm0_data_valid  ,

            // manager 27, lane 7, stream 1      
            input   wire                                        std__mgr27__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane7_strm1_data        ,
            output  wire                                        mgr27__std__lane7_strm1_data_valid  ,

            // manager 27, lane 8, stream 0      
            input   wire                                        std__mgr27__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane8_strm0_data        ,
            output  wire                                        mgr27__std__lane8_strm0_data_valid  ,

            // manager 27, lane 8, stream 1      
            input   wire                                        std__mgr27__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane8_strm1_data        ,
            output  wire                                        mgr27__std__lane8_strm1_data_valid  ,

            // manager 27, lane 9, stream 0      
            input   wire                                        std__mgr27__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane9_strm0_data        ,
            output  wire                                        mgr27__std__lane9_strm0_data_valid  ,

            // manager 27, lane 9, stream 1      
            input   wire                                        std__mgr27__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane9_strm1_data        ,
            output  wire                                        mgr27__std__lane9_strm1_data_valid  ,

            // manager 27, lane 10, stream 0      
            input   wire                                        std__mgr27__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane10_strm0_data        ,
            output  wire                                        mgr27__std__lane10_strm0_data_valid  ,

            // manager 27, lane 10, stream 1      
            input   wire                                        std__mgr27__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane10_strm1_data        ,
            output  wire                                        mgr27__std__lane10_strm1_data_valid  ,

            // manager 27, lane 11, stream 0      
            input   wire                                        std__mgr27__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane11_strm0_data        ,
            output  wire                                        mgr27__std__lane11_strm0_data_valid  ,

            // manager 27, lane 11, stream 1      
            input   wire                                        std__mgr27__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane11_strm1_data        ,
            output  wire                                        mgr27__std__lane11_strm1_data_valid  ,

            // manager 27, lane 12, stream 0      
            input   wire                                        std__mgr27__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane12_strm0_data        ,
            output  wire                                        mgr27__std__lane12_strm0_data_valid  ,

            // manager 27, lane 12, stream 1      
            input   wire                                        std__mgr27__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane12_strm1_data        ,
            output  wire                                        mgr27__std__lane12_strm1_data_valid  ,

            // manager 27, lane 13, stream 0      
            input   wire                                        std__mgr27__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane13_strm0_data        ,
            output  wire                                        mgr27__std__lane13_strm0_data_valid  ,

            // manager 27, lane 13, stream 1      
            input   wire                                        std__mgr27__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane13_strm1_data        ,
            output  wire                                        mgr27__std__lane13_strm1_data_valid  ,

            // manager 27, lane 14, stream 0      
            input   wire                                        std__mgr27__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane14_strm0_data        ,
            output  wire                                        mgr27__std__lane14_strm0_data_valid  ,

            // manager 27, lane 14, stream 1      
            input   wire                                        std__mgr27__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane14_strm1_data        ,
            output  wire                                        mgr27__std__lane14_strm1_data_valid  ,

            // manager 27, lane 15, stream 0      
            input   wire                                        std__mgr27__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane15_strm0_data        ,
            output  wire                                        mgr27__std__lane15_strm0_data_valid  ,

            // manager 27, lane 15, stream 1      
            input   wire                                        std__mgr27__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane15_strm1_data        ,
            output  wire                                        mgr27__std__lane15_strm1_data_valid  ,

            // manager 27, lane 16, stream 0      
            input   wire                                        std__mgr27__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane16_strm0_data        ,
            output  wire                                        mgr27__std__lane16_strm0_data_valid  ,

            // manager 27, lane 16, stream 1      
            input   wire                                        std__mgr27__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane16_strm1_data        ,
            output  wire                                        mgr27__std__lane16_strm1_data_valid  ,

            // manager 27, lane 17, stream 0      
            input   wire                                        std__mgr27__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane17_strm0_data        ,
            output  wire                                        mgr27__std__lane17_strm0_data_valid  ,

            // manager 27, lane 17, stream 1      
            input   wire                                        std__mgr27__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane17_strm1_data        ,
            output  wire                                        mgr27__std__lane17_strm1_data_valid  ,

            // manager 27, lane 18, stream 0      
            input   wire                                        std__mgr27__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane18_strm0_data        ,
            output  wire                                        mgr27__std__lane18_strm0_data_valid  ,

            // manager 27, lane 18, stream 1      
            input   wire                                        std__mgr27__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane18_strm1_data        ,
            output  wire                                        mgr27__std__lane18_strm1_data_valid  ,

            // manager 27, lane 19, stream 0      
            input   wire                                        std__mgr27__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane19_strm0_data        ,
            output  wire                                        mgr27__std__lane19_strm0_data_valid  ,

            // manager 27, lane 19, stream 1      
            input   wire                                        std__mgr27__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane19_strm1_data        ,
            output  wire                                        mgr27__std__lane19_strm1_data_valid  ,

            // manager 27, lane 20, stream 0      
            input   wire                                        std__mgr27__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane20_strm0_data        ,
            output  wire                                        mgr27__std__lane20_strm0_data_valid  ,

            // manager 27, lane 20, stream 1      
            input   wire                                        std__mgr27__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane20_strm1_data        ,
            output  wire                                        mgr27__std__lane20_strm1_data_valid  ,

            // manager 27, lane 21, stream 0      
            input   wire                                        std__mgr27__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane21_strm0_data        ,
            output  wire                                        mgr27__std__lane21_strm0_data_valid  ,

            // manager 27, lane 21, stream 1      
            input   wire                                        std__mgr27__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane21_strm1_data        ,
            output  wire                                        mgr27__std__lane21_strm1_data_valid  ,

            // manager 27, lane 22, stream 0      
            input   wire                                        std__mgr27__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane22_strm0_data        ,
            output  wire                                        mgr27__std__lane22_strm0_data_valid  ,

            // manager 27, lane 22, stream 1      
            input   wire                                        std__mgr27__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane22_strm1_data        ,
            output  wire                                        mgr27__std__lane22_strm1_data_valid  ,

            // manager 27, lane 23, stream 0      
            input   wire                                        std__mgr27__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane23_strm0_data        ,
            output  wire                                        mgr27__std__lane23_strm0_data_valid  ,

            // manager 27, lane 23, stream 1      
            input   wire                                        std__mgr27__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane23_strm1_data        ,
            output  wire                                        mgr27__std__lane23_strm1_data_valid  ,

            // manager 27, lane 24, stream 0      
            input   wire                                        std__mgr27__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane24_strm0_data        ,
            output  wire                                        mgr27__std__lane24_strm0_data_valid  ,

            // manager 27, lane 24, stream 1      
            input   wire                                        std__mgr27__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane24_strm1_data        ,
            output  wire                                        mgr27__std__lane24_strm1_data_valid  ,

            // manager 27, lane 25, stream 0      
            input   wire                                        std__mgr27__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane25_strm0_data        ,
            output  wire                                        mgr27__std__lane25_strm0_data_valid  ,

            // manager 27, lane 25, stream 1      
            input   wire                                        std__mgr27__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane25_strm1_data        ,
            output  wire                                        mgr27__std__lane25_strm1_data_valid  ,

            // manager 27, lane 26, stream 0      
            input   wire                                        std__mgr27__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane26_strm0_data        ,
            output  wire                                        mgr27__std__lane26_strm0_data_valid  ,

            // manager 27, lane 26, stream 1      
            input   wire                                        std__mgr27__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane26_strm1_data        ,
            output  wire                                        mgr27__std__lane26_strm1_data_valid  ,

            // manager 27, lane 27, stream 0      
            input   wire                                        std__mgr27__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane27_strm0_data        ,
            output  wire                                        mgr27__std__lane27_strm0_data_valid  ,

            // manager 27, lane 27, stream 1      
            input   wire                                        std__mgr27__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane27_strm1_data        ,
            output  wire                                        mgr27__std__lane27_strm1_data_valid  ,

            // manager 27, lane 28, stream 0      
            input   wire                                        std__mgr27__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane28_strm0_data        ,
            output  wire                                        mgr27__std__lane28_strm0_data_valid  ,

            // manager 27, lane 28, stream 1      
            input   wire                                        std__mgr27__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane28_strm1_data        ,
            output  wire                                        mgr27__std__lane28_strm1_data_valid  ,

            // manager 27, lane 29, stream 0      
            input   wire                                        std__mgr27__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane29_strm0_data        ,
            output  wire                                        mgr27__std__lane29_strm0_data_valid  ,

            // manager 27, lane 29, stream 1      
            input   wire                                        std__mgr27__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane29_strm1_data        ,
            output  wire                                        mgr27__std__lane29_strm1_data_valid  ,

            // manager 27, lane 30, stream 0      
            input   wire                                        std__mgr27__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane30_strm0_data        ,
            output  wire                                        mgr27__std__lane30_strm0_data_valid  ,

            // manager 27, lane 30, stream 1      
            input   wire                                        std__mgr27__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane30_strm1_data        ,
            output  wire                                        mgr27__std__lane30_strm1_data_valid  ,

            // manager 27, lane 31, stream 0      
            input   wire                                        std__mgr27__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane31_strm0_data        ,
            output  wire                                        mgr27__std__lane31_strm0_data_valid  ,

            // manager 27, lane 31, stream 1      
            input   wire                                        std__mgr27__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr27__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr27__std__lane31_strm1_data        ,
            output  wire                                        mgr27__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 28, lane 0, stream 0      
            input   wire                                        std__mgr28__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane0_strm0_data        ,
            output  wire                                        mgr28__std__lane0_strm0_data_valid  ,

            // manager 28, lane 0, stream 1      
            input   wire                                        std__mgr28__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane0_strm1_data        ,
            output  wire                                        mgr28__std__lane0_strm1_data_valid  ,

            // manager 28, lane 1, stream 0      
            input   wire                                        std__mgr28__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane1_strm0_data        ,
            output  wire                                        mgr28__std__lane1_strm0_data_valid  ,

            // manager 28, lane 1, stream 1      
            input   wire                                        std__mgr28__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane1_strm1_data        ,
            output  wire                                        mgr28__std__lane1_strm1_data_valid  ,

            // manager 28, lane 2, stream 0      
            input   wire                                        std__mgr28__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane2_strm0_data        ,
            output  wire                                        mgr28__std__lane2_strm0_data_valid  ,

            // manager 28, lane 2, stream 1      
            input   wire                                        std__mgr28__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane2_strm1_data        ,
            output  wire                                        mgr28__std__lane2_strm1_data_valid  ,

            // manager 28, lane 3, stream 0      
            input   wire                                        std__mgr28__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane3_strm0_data        ,
            output  wire                                        mgr28__std__lane3_strm0_data_valid  ,

            // manager 28, lane 3, stream 1      
            input   wire                                        std__mgr28__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane3_strm1_data        ,
            output  wire                                        mgr28__std__lane3_strm1_data_valid  ,

            // manager 28, lane 4, stream 0      
            input   wire                                        std__mgr28__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane4_strm0_data        ,
            output  wire                                        mgr28__std__lane4_strm0_data_valid  ,

            // manager 28, lane 4, stream 1      
            input   wire                                        std__mgr28__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane4_strm1_data        ,
            output  wire                                        mgr28__std__lane4_strm1_data_valid  ,

            // manager 28, lane 5, stream 0      
            input   wire                                        std__mgr28__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane5_strm0_data        ,
            output  wire                                        mgr28__std__lane5_strm0_data_valid  ,

            // manager 28, lane 5, stream 1      
            input   wire                                        std__mgr28__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane5_strm1_data        ,
            output  wire                                        mgr28__std__lane5_strm1_data_valid  ,

            // manager 28, lane 6, stream 0      
            input   wire                                        std__mgr28__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane6_strm0_data        ,
            output  wire                                        mgr28__std__lane6_strm0_data_valid  ,

            // manager 28, lane 6, stream 1      
            input   wire                                        std__mgr28__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane6_strm1_data        ,
            output  wire                                        mgr28__std__lane6_strm1_data_valid  ,

            // manager 28, lane 7, stream 0      
            input   wire                                        std__mgr28__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane7_strm0_data        ,
            output  wire                                        mgr28__std__lane7_strm0_data_valid  ,

            // manager 28, lane 7, stream 1      
            input   wire                                        std__mgr28__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane7_strm1_data        ,
            output  wire                                        mgr28__std__lane7_strm1_data_valid  ,

            // manager 28, lane 8, stream 0      
            input   wire                                        std__mgr28__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane8_strm0_data        ,
            output  wire                                        mgr28__std__lane8_strm0_data_valid  ,

            // manager 28, lane 8, stream 1      
            input   wire                                        std__mgr28__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane8_strm1_data        ,
            output  wire                                        mgr28__std__lane8_strm1_data_valid  ,

            // manager 28, lane 9, stream 0      
            input   wire                                        std__mgr28__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane9_strm0_data        ,
            output  wire                                        mgr28__std__lane9_strm0_data_valid  ,

            // manager 28, lane 9, stream 1      
            input   wire                                        std__mgr28__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane9_strm1_data        ,
            output  wire                                        mgr28__std__lane9_strm1_data_valid  ,

            // manager 28, lane 10, stream 0      
            input   wire                                        std__mgr28__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane10_strm0_data        ,
            output  wire                                        mgr28__std__lane10_strm0_data_valid  ,

            // manager 28, lane 10, stream 1      
            input   wire                                        std__mgr28__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane10_strm1_data        ,
            output  wire                                        mgr28__std__lane10_strm1_data_valid  ,

            // manager 28, lane 11, stream 0      
            input   wire                                        std__mgr28__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane11_strm0_data        ,
            output  wire                                        mgr28__std__lane11_strm0_data_valid  ,

            // manager 28, lane 11, stream 1      
            input   wire                                        std__mgr28__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane11_strm1_data        ,
            output  wire                                        mgr28__std__lane11_strm1_data_valid  ,

            // manager 28, lane 12, stream 0      
            input   wire                                        std__mgr28__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane12_strm0_data        ,
            output  wire                                        mgr28__std__lane12_strm0_data_valid  ,

            // manager 28, lane 12, stream 1      
            input   wire                                        std__mgr28__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane12_strm1_data        ,
            output  wire                                        mgr28__std__lane12_strm1_data_valid  ,

            // manager 28, lane 13, stream 0      
            input   wire                                        std__mgr28__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane13_strm0_data        ,
            output  wire                                        mgr28__std__lane13_strm0_data_valid  ,

            // manager 28, lane 13, stream 1      
            input   wire                                        std__mgr28__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane13_strm1_data        ,
            output  wire                                        mgr28__std__lane13_strm1_data_valid  ,

            // manager 28, lane 14, stream 0      
            input   wire                                        std__mgr28__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane14_strm0_data        ,
            output  wire                                        mgr28__std__lane14_strm0_data_valid  ,

            // manager 28, lane 14, stream 1      
            input   wire                                        std__mgr28__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane14_strm1_data        ,
            output  wire                                        mgr28__std__lane14_strm1_data_valid  ,

            // manager 28, lane 15, stream 0      
            input   wire                                        std__mgr28__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane15_strm0_data        ,
            output  wire                                        mgr28__std__lane15_strm0_data_valid  ,

            // manager 28, lane 15, stream 1      
            input   wire                                        std__mgr28__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane15_strm1_data        ,
            output  wire                                        mgr28__std__lane15_strm1_data_valid  ,

            // manager 28, lane 16, stream 0      
            input   wire                                        std__mgr28__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane16_strm0_data        ,
            output  wire                                        mgr28__std__lane16_strm0_data_valid  ,

            // manager 28, lane 16, stream 1      
            input   wire                                        std__mgr28__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane16_strm1_data        ,
            output  wire                                        mgr28__std__lane16_strm1_data_valid  ,

            // manager 28, lane 17, stream 0      
            input   wire                                        std__mgr28__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane17_strm0_data        ,
            output  wire                                        mgr28__std__lane17_strm0_data_valid  ,

            // manager 28, lane 17, stream 1      
            input   wire                                        std__mgr28__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane17_strm1_data        ,
            output  wire                                        mgr28__std__lane17_strm1_data_valid  ,

            // manager 28, lane 18, stream 0      
            input   wire                                        std__mgr28__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane18_strm0_data        ,
            output  wire                                        mgr28__std__lane18_strm0_data_valid  ,

            // manager 28, lane 18, stream 1      
            input   wire                                        std__mgr28__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane18_strm1_data        ,
            output  wire                                        mgr28__std__lane18_strm1_data_valid  ,

            // manager 28, lane 19, stream 0      
            input   wire                                        std__mgr28__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane19_strm0_data        ,
            output  wire                                        mgr28__std__lane19_strm0_data_valid  ,

            // manager 28, lane 19, stream 1      
            input   wire                                        std__mgr28__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane19_strm1_data        ,
            output  wire                                        mgr28__std__lane19_strm1_data_valid  ,

            // manager 28, lane 20, stream 0      
            input   wire                                        std__mgr28__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane20_strm0_data        ,
            output  wire                                        mgr28__std__lane20_strm0_data_valid  ,

            // manager 28, lane 20, stream 1      
            input   wire                                        std__mgr28__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane20_strm1_data        ,
            output  wire                                        mgr28__std__lane20_strm1_data_valid  ,

            // manager 28, lane 21, stream 0      
            input   wire                                        std__mgr28__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane21_strm0_data        ,
            output  wire                                        mgr28__std__lane21_strm0_data_valid  ,

            // manager 28, lane 21, stream 1      
            input   wire                                        std__mgr28__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane21_strm1_data        ,
            output  wire                                        mgr28__std__lane21_strm1_data_valid  ,

            // manager 28, lane 22, stream 0      
            input   wire                                        std__mgr28__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane22_strm0_data        ,
            output  wire                                        mgr28__std__lane22_strm0_data_valid  ,

            // manager 28, lane 22, stream 1      
            input   wire                                        std__mgr28__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane22_strm1_data        ,
            output  wire                                        mgr28__std__lane22_strm1_data_valid  ,

            // manager 28, lane 23, stream 0      
            input   wire                                        std__mgr28__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane23_strm0_data        ,
            output  wire                                        mgr28__std__lane23_strm0_data_valid  ,

            // manager 28, lane 23, stream 1      
            input   wire                                        std__mgr28__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane23_strm1_data        ,
            output  wire                                        mgr28__std__lane23_strm1_data_valid  ,

            // manager 28, lane 24, stream 0      
            input   wire                                        std__mgr28__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane24_strm0_data        ,
            output  wire                                        mgr28__std__lane24_strm0_data_valid  ,

            // manager 28, lane 24, stream 1      
            input   wire                                        std__mgr28__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane24_strm1_data        ,
            output  wire                                        mgr28__std__lane24_strm1_data_valid  ,

            // manager 28, lane 25, stream 0      
            input   wire                                        std__mgr28__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane25_strm0_data        ,
            output  wire                                        mgr28__std__lane25_strm0_data_valid  ,

            // manager 28, lane 25, stream 1      
            input   wire                                        std__mgr28__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane25_strm1_data        ,
            output  wire                                        mgr28__std__lane25_strm1_data_valid  ,

            // manager 28, lane 26, stream 0      
            input   wire                                        std__mgr28__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane26_strm0_data        ,
            output  wire                                        mgr28__std__lane26_strm0_data_valid  ,

            // manager 28, lane 26, stream 1      
            input   wire                                        std__mgr28__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane26_strm1_data        ,
            output  wire                                        mgr28__std__lane26_strm1_data_valid  ,

            // manager 28, lane 27, stream 0      
            input   wire                                        std__mgr28__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane27_strm0_data        ,
            output  wire                                        mgr28__std__lane27_strm0_data_valid  ,

            // manager 28, lane 27, stream 1      
            input   wire                                        std__mgr28__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane27_strm1_data        ,
            output  wire                                        mgr28__std__lane27_strm1_data_valid  ,

            // manager 28, lane 28, stream 0      
            input   wire                                        std__mgr28__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane28_strm0_data        ,
            output  wire                                        mgr28__std__lane28_strm0_data_valid  ,

            // manager 28, lane 28, stream 1      
            input   wire                                        std__mgr28__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane28_strm1_data        ,
            output  wire                                        mgr28__std__lane28_strm1_data_valid  ,

            // manager 28, lane 29, stream 0      
            input   wire                                        std__mgr28__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane29_strm0_data        ,
            output  wire                                        mgr28__std__lane29_strm0_data_valid  ,

            // manager 28, lane 29, stream 1      
            input   wire                                        std__mgr28__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane29_strm1_data        ,
            output  wire                                        mgr28__std__lane29_strm1_data_valid  ,

            // manager 28, lane 30, stream 0      
            input   wire                                        std__mgr28__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane30_strm0_data        ,
            output  wire                                        mgr28__std__lane30_strm0_data_valid  ,

            // manager 28, lane 30, stream 1      
            input   wire                                        std__mgr28__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane30_strm1_data        ,
            output  wire                                        mgr28__std__lane30_strm1_data_valid  ,

            // manager 28, lane 31, stream 0      
            input   wire                                        std__mgr28__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane31_strm0_data        ,
            output  wire                                        mgr28__std__lane31_strm0_data_valid  ,

            // manager 28, lane 31, stream 1      
            input   wire                                        std__mgr28__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr28__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr28__std__lane31_strm1_data        ,
            output  wire                                        mgr28__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 29, lane 0, stream 0      
            input   wire                                        std__mgr29__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane0_strm0_data        ,
            output  wire                                        mgr29__std__lane0_strm0_data_valid  ,

            // manager 29, lane 0, stream 1      
            input   wire                                        std__mgr29__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane0_strm1_data        ,
            output  wire                                        mgr29__std__lane0_strm1_data_valid  ,

            // manager 29, lane 1, stream 0      
            input   wire                                        std__mgr29__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane1_strm0_data        ,
            output  wire                                        mgr29__std__lane1_strm0_data_valid  ,

            // manager 29, lane 1, stream 1      
            input   wire                                        std__mgr29__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane1_strm1_data        ,
            output  wire                                        mgr29__std__lane1_strm1_data_valid  ,

            // manager 29, lane 2, stream 0      
            input   wire                                        std__mgr29__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane2_strm0_data        ,
            output  wire                                        mgr29__std__lane2_strm0_data_valid  ,

            // manager 29, lane 2, stream 1      
            input   wire                                        std__mgr29__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane2_strm1_data        ,
            output  wire                                        mgr29__std__lane2_strm1_data_valid  ,

            // manager 29, lane 3, stream 0      
            input   wire                                        std__mgr29__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane3_strm0_data        ,
            output  wire                                        mgr29__std__lane3_strm0_data_valid  ,

            // manager 29, lane 3, stream 1      
            input   wire                                        std__mgr29__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane3_strm1_data        ,
            output  wire                                        mgr29__std__lane3_strm1_data_valid  ,

            // manager 29, lane 4, stream 0      
            input   wire                                        std__mgr29__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane4_strm0_data        ,
            output  wire                                        mgr29__std__lane4_strm0_data_valid  ,

            // manager 29, lane 4, stream 1      
            input   wire                                        std__mgr29__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane4_strm1_data        ,
            output  wire                                        mgr29__std__lane4_strm1_data_valid  ,

            // manager 29, lane 5, stream 0      
            input   wire                                        std__mgr29__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane5_strm0_data        ,
            output  wire                                        mgr29__std__lane5_strm0_data_valid  ,

            // manager 29, lane 5, stream 1      
            input   wire                                        std__mgr29__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane5_strm1_data        ,
            output  wire                                        mgr29__std__lane5_strm1_data_valid  ,

            // manager 29, lane 6, stream 0      
            input   wire                                        std__mgr29__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane6_strm0_data        ,
            output  wire                                        mgr29__std__lane6_strm0_data_valid  ,

            // manager 29, lane 6, stream 1      
            input   wire                                        std__mgr29__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane6_strm1_data        ,
            output  wire                                        mgr29__std__lane6_strm1_data_valid  ,

            // manager 29, lane 7, stream 0      
            input   wire                                        std__mgr29__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane7_strm0_data        ,
            output  wire                                        mgr29__std__lane7_strm0_data_valid  ,

            // manager 29, lane 7, stream 1      
            input   wire                                        std__mgr29__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane7_strm1_data        ,
            output  wire                                        mgr29__std__lane7_strm1_data_valid  ,

            // manager 29, lane 8, stream 0      
            input   wire                                        std__mgr29__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane8_strm0_data        ,
            output  wire                                        mgr29__std__lane8_strm0_data_valid  ,

            // manager 29, lane 8, stream 1      
            input   wire                                        std__mgr29__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane8_strm1_data        ,
            output  wire                                        mgr29__std__lane8_strm1_data_valid  ,

            // manager 29, lane 9, stream 0      
            input   wire                                        std__mgr29__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane9_strm0_data        ,
            output  wire                                        mgr29__std__lane9_strm0_data_valid  ,

            // manager 29, lane 9, stream 1      
            input   wire                                        std__mgr29__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane9_strm1_data        ,
            output  wire                                        mgr29__std__lane9_strm1_data_valid  ,

            // manager 29, lane 10, stream 0      
            input   wire                                        std__mgr29__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane10_strm0_data        ,
            output  wire                                        mgr29__std__lane10_strm0_data_valid  ,

            // manager 29, lane 10, stream 1      
            input   wire                                        std__mgr29__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane10_strm1_data        ,
            output  wire                                        mgr29__std__lane10_strm1_data_valid  ,

            // manager 29, lane 11, stream 0      
            input   wire                                        std__mgr29__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane11_strm0_data        ,
            output  wire                                        mgr29__std__lane11_strm0_data_valid  ,

            // manager 29, lane 11, stream 1      
            input   wire                                        std__mgr29__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane11_strm1_data        ,
            output  wire                                        mgr29__std__lane11_strm1_data_valid  ,

            // manager 29, lane 12, stream 0      
            input   wire                                        std__mgr29__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane12_strm0_data        ,
            output  wire                                        mgr29__std__lane12_strm0_data_valid  ,

            // manager 29, lane 12, stream 1      
            input   wire                                        std__mgr29__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane12_strm1_data        ,
            output  wire                                        mgr29__std__lane12_strm1_data_valid  ,

            // manager 29, lane 13, stream 0      
            input   wire                                        std__mgr29__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane13_strm0_data        ,
            output  wire                                        mgr29__std__lane13_strm0_data_valid  ,

            // manager 29, lane 13, stream 1      
            input   wire                                        std__mgr29__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane13_strm1_data        ,
            output  wire                                        mgr29__std__lane13_strm1_data_valid  ,

            // manager 29, lane 14, stream 0      
            input   wire                                        std__mgr29__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane14_strm0_data        ,
            output  wire                                        mgr29__std__lane14_strm0_data_valid  ,

            // manager 29, lane 14, stream 1      
            input   wire                                        std__mgr29__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane14_strm1_data        ,
            output  wire                                        mgr29__std__lane14_strm1_data_valid  ,

            // manager 29, lane 15, stream 0      
            input   wire                                        std__mgr29__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane15_strm0_data        ,
            output  wire                                        mgr29__std__lane15_strm0_data_valid  ,

            // manager 29, lane 15, stream 1      
            input   wire                                        std__mgr29__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane15_strm1_data        ,
            output  wire                                        mgr29__std__lane15_strm1_data_valid  ,

            // manager 29, lane 16, stream 0      
            input   wire                                        std__mgr29__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane16_strm0_data        ,
            output  wire                                        mgr29__std__lane16_strm0_data_valid  ,

            // manager 29, lane 16, stream 1      
            input   wire                                        std__mgr29__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane16_strm1_data        ,
            output  wire                                        mgr29__std__lane16_strm1_data_valid  ,

            // manager 29, lane 17, stream 0      
            input   wire                                        std__mgr29__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane17_strm0_data        ,
            output  wire                                        mgr29__std__lane17_strm0_data_valid  ,

            // manager 29, lane 17, stream 1      
            input   wire                                        std__mgr29__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane17_strm1_data        ,
            output  wire                                        mgr29__std__lane17_strm1_data_valid  ,

            // manager 29, lane 18, stream 0      
            input   wire                                        std__mgr29__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane18_strm0_data        ,
            output  wire                                        mgr29__std__lane18_strm0_data_valid  ,

            // manager 29, lane 18, stream 1      
            input   wire                                        std__mgr29__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane18_strm1_data        ,
            output  wire                                        mgr29__std__lane18_strm1_data_valid  ,

            // manager 29, lane 19, stream 0      
            input   wire                                        std__mgr29__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane19_strm0_data        ,
            output  wire                                        mgr29__std__lane19_strm0_data_valid  ,

            // manager 29, lane 19, stream 1      
            input   wire                                        std__mgr29__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane19_strm1_data        ,
            output  wire                                        mgr29__std__lane19_strm1_data_valid  ,

            // manager 29, lane 20, stream 0      
            input   wire                                        std__mgr29__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane20_strm0_data        ,
            output  wire                                        mgr29__std__lane20_strm0_data_valid  ,

            // manager 29, lane 20, stream 1      
            input   wire                                        std__mgr29__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane20_strm1_data        ,
            output  wire                                        mgr29__std__lane20_strm1_data_valid  ,

            // manager 29, lane 21, stream 0      
            input   wire                                        std__mgr29__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane21_strm0_data        ,
            output  wire                                        mgr29__std__lane21_strm0_data_valid  ,

            // manager 29, lane 21, stream 1      
            input   wire                                        std__mgr29__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane21_strm1_data        ,
            output  wire                                        mgr29__std__lane21_strm1_data_valid  ,

            // manager 29, lane 22, stream 0      
            input   wire                                        std__mgr29__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane22_strm0_data        ,
            output  wire                                        mgr29__std__lane22_strm0_data_valid  ,

            // manager 29, lane 22, stream 1      
            input   wire                                        std__mgr29__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane22_strm1_data        ,
            output  wire                                        mgr29__std__lane22_strm1_data_valid  ,

            // manager 29, lane 23, stream 0      
            input   wire                                        std__mgr29__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane23_strm0_data        ,
            output  wire                                        mgr29__std__lane23_strm0_data_valid  ,

            // manager 29, lane 23, stream 1      
            input   wire                                        std__mgr29__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane23_strm1_data        ,
            output  wire                                        mgr29__std__lane23_strm1_data_valid  ,

            // manager 29, lane 24, stream 0      
            input   wire                                        std__mgr29__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane24_strm0_data        ,
            output  wire                                        mgr29__std__lane24_strm0_data_valid  ,

            // manager 29, lane 24, stream 1      
            input   wire                                        std__mgr29__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane24_strm1_data        ,
            output  wire                                        mgr29__std__lane24_strm1_data_valid  ,

            // manager 29, lane 25, stream 0      
            input   wire                                        std__mgr29__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane25_strm0_data        ,
            output  wire                                        mgr29__std__lane25_strm0_data_valid  ,

            // manager 29, lane 25, stream 1      
            input   wire                                        std__mgr29__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane25_strm1_data        ,
            output  wire                                        mgr29__std__lane25_strm1_data_valid  ,

            // manager 29, lane 26, stream 0      
            input   wire                                        std__mgr29__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane26_strm0_data        ,
            output  wire                                        mgr29__std__lane26_strm0_data_valid  ,

            // manager 29, lane 26, stream 1      
            input   wire                                        std__mgr29__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane26_strm1_data        ,
            output  wire                                        mgr29__std__lane26_strm1_data_valid  ,

            // manager 29, lane 27, stream 0      
            input   wire                                        std__mgr29__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane27_strm0_data        ,
            output  wire                                        mgr29__std__lane27_strm0_data_valid  ,

            // manager 29, lane 27, stream 1      
            input   wire                                        std__mgr29__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane27_strm1_data        ,
            output  wire                                        mgr29__std__lane27_strm1_data_valid  ,

            // manager 29, lane 28, stream 0      
            input   wire                                        std__mgr29__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane28_strm0_data        ,
            output  wire                                        mgr29__std__lane28_strm0_data_valid  ,

            // manager 29, lane 28, stream 1      
            input   wire                                        std__mgr29__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane28_strm1_data        ,
            output  wire                                        mgr29__std__lane28_strm1_data_valid  ,

            // manager 29, lane 29, stream 0      
            input   wire                                        std__mgr29__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane29_strm0_data        ,
            output  wire                                        mgr29__std__lane29_strm0_data_valid  ,

            // manager 29, lane 29, stream 1      
            input   wire                                        std__mgr29__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane29_strm1_data        ,
            output  wire                                        mgr29__std__lane29_strm1_data_valid  ,

            // manager 29, lane 30, stream 0      
            input   wire                                        std__mgr29__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane30_strm0_data        ,
            output  wire                                        mgr29__std__lane30_strm0_data_valid  ,

            // manager 29, lane 30, stream 1      
            input   wire                                        std__mgr29__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane30_strm1_data        ,
            output  wire                                        mgr29__std__lane30_strm1_data_valid  ,

            // manager 29, lane 31, stream 0      
            input   wire                                        std__mgr29__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane31_strm0_data        ,
            output  wire                                        mgr29__std__lane31_strm0_data_valid  ,

            // manager 29, lane 31, stream 1      
            input   wire                                        std__mgr29__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr29__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr29__std__lane31_strm1_data        ,
            output  wire                                        mgr29__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 30, lane 0, stream 0      
            input   wire                                        std__mgr30__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane0_strm0_data        ,
            output  wire                                        mgr30__std__lane0_strm0_data_valid  ,

            // manager 30, lane 0, stream 1      
            input   wire                                        std__mgr30__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane0_strm1_data        ,
            output  wire                                        mgr30__std__lane0_strm1_data_valid  ,

            // manager 30, lane 1, stream 0      
            input   wire                                        std__mgr30__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane1_strm0_data        ,
            output  wire                                        mgr30__std__lane1_strm0_data_valid  ,

            // manager 30, lane 1, stream 1      
            input   wire                                        std__mgr30__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane1_strm1_data        ,
            output  wire                                        mgr30__std__lane1_strm1_data_valid  ,

            // manager 30, lane 2, stream 0      
            input   wire                                        std__mgr30__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane2_strm0_data        ,
            output  wire                                        mgr30__std__lane2_strm0_data_valid  ,

            // manager 30, lane 2, stream 1      
            input   wire                                        std__mgr30__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane2_strm1_data        ,
            output  wire                                        mgr30__std__lane2_strm1_data_valid  ,

            // manager 30, lane 3, stream 0      
            input   wire                                        std__mgr30__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane3_strm0_data        ,
            output  wire                                        mgr30__std__lane3_strm0_data_valid  ,

            // manager 30, lane 3, stream 1      
            input   wire                                        std__mgr30__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane3_strm1_data        ,
            output  wire                                        mgr30__std__lane3_strm1_data_valid  ,

            // manager 30, lane 4, stream 0      
            input   wire                                        std__mgr30__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane4_strm0_data        ,
            output  wire                                        mgr30__std__lane4_strm0_data_valid  ,

            // manager 30, lane 4, stream 1      
            input   wire                                        std__mgr30__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane4_strm1_data        ,
            output  wire                                        mgr30__std__lane4_strm1_data_valid  ,

            // manager 30, lane 5, stream 0      
            input   wire                                        std__mgr30__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane5_strm0_data        ,
            output  wire                                        mgr30__std__lane5_strm0_data_valid  ,

            // manager 30, lane 5, stream 1      
            input   wire                                        std__mgr30__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane5_strm1_data        ,
            output  wire                                        mgr30__std__lane5_strm1_data_valid  ,

            // manager 30, lane 6, stream 0      
            input   wire                                        std__mgr30__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane6_strm0_data        ,
            output  wire                                        mgr30__std__lane6_strm0_data_valid  ,

            // manager 30, lane 6, stream 1      
            input   wire                                        std__mgr30__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane6_strm1_data        ,
            output  wire                                        mgr30__std__lane6_strm1_data_valid  ,

            // manager 30, lane 7, stream 0      
            input   wire                                        std__mgr30__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane7_strm0_data        ,
            output  wire                                        mgr30__std__lane7_strm0_data_valid  ,

            // manager 30, lane 7, stream 1      
            input   wire                                        std__mgr30__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane7_strm1_data        ,
            output  wire                                        mgr30__std__lane7_strm1_data_valid  ,

            // manager 30, lane 8, stream 0      
            input   wire                                        std__mgr30__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane8_strm0_data        ,
            output  wire                                        mgr30__std__lane8_strm0_data_valid  ,

            // manager 30, lane 8, stream 1      
            input   wire                                        std__mgr30__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane8_strm1_data        ,
            output  wire                                        mgr30__std__lane8_strm1_data_valid  ,

            // manager 30, lane 9, stream 0      
            input   wire                                        std__mgr30__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane9_strm0_data        ,
            output  wire                                        mgr30__std__lane9_strm0_data_valid  ,

            // manager 30, lane 9, stream 1      
            input   wire                                        std__mgr30__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane9_strm1_data        ,
            output  wire                                        mgr30__std__lane9_strm1_data_valid  ,

            // manager 30, lane 10, stream 0      
            input   wire                                        std__mgr30__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane10_strm0_data        ,
            output  wire                                        mgr30__std__lane10_strm0_data_valid  ,

            // manager 30, lane 10, stream 1      
            input   wire                                        std__mgr30__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane10_strm1_data        ,
            output  wire                                        mgr30__std__lane10_strm1_data_valid  ,

            // manager 30, lane 11, stream 0      
            input   wire                                        std__mgr30__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane11_strm0_data        ,
            output  wire                                        mgr30__std__lane11_strm0_data_valid  ,

            // manager 30, lane 11, stream 1      
            input   wire                                        std__mgr30__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane11_strm1_data        ,
            output  wire                                        mgr30__std__lane11_strm1_data_valid  ,

            // manager 30, lane 12, stream 0      
            input   wire                                        std__mgr30__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane12_strm0_data        ,
            output  wire                                        mgr30__std__lane12_strm0_data_valid  ,

            // manager 30, lane 12, stream 1      
            input   wire                                        std__mgr30__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane12_strm1_data        ,
            output  wire                                        mgr30__std__lane12_strm1_data_valid  ,

            // manager 30, lane 13, stream 0      
            input   wire                                        std__mgr30__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane13_strm0_data        ,
            output  wire                                        mgr30__std__lane13_strm0_data_valid  ,

            // manager 30, lane 13, stream 1      
            input   wire                                        std__mgr30__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane13_strm1_data        ,
            output  wire                                        mgr30__std__lane13_strm1_data_valid  ,

            // manager 30, lane 14, stream 0      
            input   wire                                        std__mgr30__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane14_strm0_data        ,
            output  wire                                        mgr30__std__lane14_strm0_data_valid  ,

            // manager 30, lane 14, stream 1      
            input   wire                                        std__mgr30__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane14_strm1_data        ,
            output  wire                                        mgr30__std__lane14_strm1_data_valid  ,

            // manager 30, lane 15, stream 0      
            input   wire                                        std__mgr30__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane15_strm0_data        ,
            output  wire                                        mgr30__std__lane15_strm0_data_valid  ,

            // manager 30, lane 15, stream 1      
            input   wire                                        std__mgr30__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane15_strm1_data        ,
            output  wire                                        mgr30__std__lane15_strm1_data_valid  ,

            // manager 30, lane 16, stream 0      
            input   wire                                        std__mgr30__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane16_strm0_data        ,
            output  wire                                        mgr30__std__lane16_strm0_data_valid  ,

            // manager 30, lane 16, stream 1      
            input   wire                                        std__mgr30__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane16_strm1_data        ,
            output  wire                                        mgr30__std__lane16_strm1_data_valid  ,

            // manager 30, lane 17, stream 0      
            input   wire                                        std__mgr30__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane17_strm0_data        ,
            output  wire                                        mgr30__std__lane17_strm0_data_valid  ,

            // manager 30, lane 17, stream 1      
            input   wire                                        std__mgr30__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane17_strm1_data        ,
            output  wire                                        mgr30__std__lane17_strm1_data_valid  ,

            // manager 30, lane 18, stream 0      
            input   wire                                        std__mgr30__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane18_strm0_data        ,
            output  wire                                        mgr30__std__lane18_strm0_data_valid  ,

            // manager 30, lane 18, stream 1      
            input   wire                                        std__mgr30__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane18_strm1_data        ,
            output  wire                                        mgr30__std__lane18_strm1_data_valid  ,

            // manager 30, lane 19, stream 0      
            input   wire                                        std__mgr30__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane19_strm0_data        ,
            output  wire                                        mgr30__std__lane19_strm0_data_valid  ,

            // manager 30, lane 19, stream 1      
            input   wire                                        std__mgr30__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane19_strm1_data        ,
            output  wire                                        mgr30__std__lane19_strm1_data_valid  ,

            // manager 30, lane 20, stream 0      
            input   wire                                        std__mgr30__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane20_strm0_data        ,
            output  wire                                        mgr30__std__lane20_strm0_data_valid  ,

            // manager 30, lane 20, stream 1      
            input   wire                                        std__mgr30__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane20_strm1_data        ,
            output  wire                                        mgr30__std__lane20_strm1_data_valid  ,

            // manager 30, lane 21, stream 0      
            input   wire                                        std__mgr30__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane21_strm0_data        ,
            output  wire                                        mgr30__std__lane21_strm0_data_valid  ,

            // manager 30, lane 21, stream 1      
            input   wire                                        std__mgr30__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane21_strm1_data        ,
            output  wire                                        mgr30__std__lane21_strm1_data_valid  ,

            // manager 30, lane 22, stream 0      
            input   wire                                        std__mgr30__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane22_strm0_data        ,
            output  wire                                        mgr30__std__lane22_strm0_data_valid  ,

            // manager 30, lane 22, stream 1      
            input   wire                                        std__mgr30__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane22_strm1_data        ,
            output  wire                                        mgr30__std__lane22_strm1_data_valid  ,

            // manager 30, lane 23, stream 0      
            input   wire                                        std__mgr30__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane23_strm0_data        ,
            output  wire                                        mgr30__std__lane23_strm0_data_valid  ,

            // manager 30, lane 23, stream 1      
            input   wire                                        std__mgr30__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane23_strm1_data        ,
            output  wire                                        mgr30__std__lane23_strm1_data_valid  ,

            // manager 30, lane 24, stream 0      
            input   wire                                        std__mgr30__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane24_strm0_data        ,
            output  wire                                        mgr30__std__lane24_strm0_data_valid  ,

            // manager 30, lane 24, stream 1      
            input   wire                                        std__mgr30__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane24_strm1_data        ,
            output  wire                                        mgr30__std__lane24_strm1_data_valid  ,

            // manager 30, lane 25, stream 0      
            input   wire                                        std__mgr30__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane25_strm0_data        ,
            output  wire                                        mgr30__std__lane25_strm0_data_valid  ,

            // manager 30, lane 25, stream 1      
            input   wire                                        std__mgr30__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane25_strm1_data        ,
            output  wire                                        mgr30__std__lane25_strm1_data_valid  ,

            // manager 30, lane 26, stream 0      
            input   wire                                        std__mgr30__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane26_strm0_data        ,
            output  wire                                        mgr30__std__lane26_strm0_data_valid  ,

            // manager 30, lane 26, stream 1      
            input   wire                                        std__mgr30__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane26_strm1_data        ,
            output  wire                                        mgr30__std__lane26_strm1_data_valid  ,

            // manager 30, lane 27, stream 0      
            input   wire                                        std__mgr30__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane27_strm0_data        ,
            output  wire                                        mgr30__std__lane27_strm0_data_valid  ,

            // manager 30, lane 27, stream 1      
            input   wire                                        std__mgr30__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane27_strm1_data        ,
            output  wire                                        mgr30__std__lane27_strm1_data_valid  ,

            // manager 30, lane 28, stream 0      
            input   wire                                        std__mgr30__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane28_strm0_data        ,
            output  wire                                        mgr30__std__lane28_strm0_data_valid  ,

            // manager 30, lane 28, stream 1      
            input   wire                                        std__mgr30__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane28_strm1_data        ,
            output  wire                                        mgr30__std__lane28_strm1_data_valid  ,

            // manager 30, lane 29, stream 0      
            input   wire                                        std__mgr30__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane29_strm0_data        ,
            output  wire                                        mgr30__std__lane29_strm0_data_valid  ,

            // manager 30, lane 29, stream 1      
            input   wire                                        std__mgr30__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane29_strm1_data        ,
            output  wire                                        mgr30__std__lane29_strm1_data_valid  ,

            // manager 30, lane 30, stream 0      
            input   wire                                        std__mgr30__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane30_strm0_data        ,
            output  wire                                        mgr30__std__lane30_strm0_data_valid  ,

            // manager 30, lane 30, stream 1      
            input   wire                                        std__mgr30__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane30_strm1_data        ,
            output  wire                                        mgr30__std__lane30_strm1_data_valid  ,

            // manager 30, lane 31, stream 0      
            input   wire                                        std__mgr30__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane31_strm0_data        ,
            output  wire                                        mgr30__std__lane31_strm0_data_valid  ,

            // manager 30, lane 31, stream 1      
            input   wire                                        std__mgr30__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr30__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr30__std__lane31_strm1_data        ,
            output  wire                                        mgr30__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 31, lane 0, stream 0      
            input   wire                                        std__mgr31__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane0_strm0_data        ,
            output  wire                                        mgr31__std__lane0_strm0_data_valid  ,

            // manager 31, lane 0, stream 1      
            input   wire                                        std__mgr31__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane0_strm1_data        ,
            output  wire                                        mgr31__std__lane0_strm1_data_valid  ,

            // manager 31, lane 1, stream 0      
            input   wire                                        std__mgr31__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane1_strm0_data        ,
            output  wire                                        mgr31__std__lane1_strm0_data_valid  ,

            // manager 31, lane 1, stream 1      
            input   wire                                        std__mgr31__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane1_strm1_data        ,
            output  wire                                        mgr31__std__lane1_strm1_data_valid  ,

            // manager 31, lane 2, stream 0      
            input   wire                                        std__mgr31__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane2_strm0_data        ,
            output  wire                                        mgr31__std__lane2_strm0_data_valid  ,

            // manager 31, lane 2, stream 1      
            input   wire                                        std__mgr31__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane2_strm1_data        ,
            output  wire                                        mgr31__std__lane2_strm1_data_valid  ,

            // manager 31, lane 3, stream 0      
            input   wire                                        std__mgr31__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane3_strm0_data        ,
            output  wire                                        mgr31__std__lane3_strm0_data_valid  ,

            // manager 31, lane 3, stream 1      
            input   wire                                        std__mgr31__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane3_strm1_data        ,
            output  wire                                        mgr31__std__lane3_strm1_data_valid  ,

            // manager 31, lane 4, stream 0      
            input   wire                                        std__mgr31__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane4_strm0_data        ,
            output  wire                                        mgr31__std__lane4_strm0_data_valid  ,

            // manager 31, lane 4, stream 1      
            input   wire                                        std__mgr31__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane4_strm1_data        ,
            output  wire                                        mgr31__std__lane4_strm1_data_valid  ,

            // manager 31, lane 5, stream 0      
            input   wire                                        std__mgr31__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane5_strm0_data        ,
            output  wire                                        mgr31__std__lane5_strm0_data_valid  ,

            // manager 31, lane 5, stream 1      
            input   wire                                        std__mgr31__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane5_strm1_data        ,
            output  wire                                        mgr31__std__lane5_strm1_data_valid  ,

            // manager 31, lane 6, stream 0      
            input   wire                                        std__mgr31__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane6_strm0_data        ,
            output  wire                                        mgr31__std__lane6_strm0_data_valid  ,

            // manager 31, lane 6, stream 1      
            input   wire                                        std__mgr31__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane6_strm1_data        ,
            output  wire                                        mgr31__std__lane6_strm1_data_valid  ,

            // manager 31, lane 7, stream 0      
            input   wire                                        std__mgr31__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane7_strm0_data        ,
            output  wire                                        mgr31__std__lane7_strm0_data_valid  ,

            // manager 31, lane 7, stream 1      
            input   wire                                        std__mgr31__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane7_strm1_data        ,
            output  wire                                        mgr31__std__lane7_strm1_data_valid  ,

            // manager 31, lane 8, stream 0      
            input   wire                                        std__mgr31__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane8_strm0_data        ,
            output  wire                                        mgr31__std__lane8_strm0_data_valid  ,

            // manager 31, lane 8, stream 1      
            input   wire                                        std__mgr31__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane8_strm1_data        ,
            output  wire                                        mgr31__std__lane8_strm1_data_valid  ,

            // manager 31, lane 9, stream 0      
            input   wire                                        std__mgr31__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane9_strm0_data        ,
            output  wire                                        mgr31__std__lane9_strm0_data_valid  ,

            // manager 31, lane 9, stream 1      
            input   wire                                        std__mgr31__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane9_strm1_data        ,
            output  wire                                        mgr31__std__lane9_strm1_data_valid  ,

            // manager 31, lane 10, stream 0      
            input   wire                                        std__mgr31__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane10_strm0_data        ,
            output  wire                                        mgr31__std__lane10_strm0_data_valid  ,

            // manager 31, lane 10, stream 1      
            input   wire                                        std__mgr31__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane10_strm1_data        ,
            output  wire                                        mgr31__std__lane10_strm1_data_valid  ,

            // manager 31, lane 11, stream 0      
            input   wire                                        std__mgr31__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane11_strm0_data        ,
            output  wire                                        mgr31__std__lane11_strm0_data_valid  ,

            // manager 31, lane 11, stream 1      
            input   wire                                        std__mgr31__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane11_strm1_data        ,
            output  wire                                        mgr31__std__lane11_strm1_data_valid  ,

            // manager 31, lane 12, stream 0      
            input   wire                                        std__mgr31__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane12_strm0_data        ,
            output  wire                                        mgr31__std__lane12_strm0_data_valid  ,

            // manager 31, lane 12, stream 1      
            input   wire                                        std__mgr31__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane12_strm1_data        ,
            output  wire                                        mgr31__std__lane12_strm1_data_valid  ,

            // manager 31, lane 13, stream 0      
            input   wire                                        std__mgr31__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane13_strm0_data        ,
            output  wire                                        mgr31__std__lane13_strm0_data_valid  ,

            // manager 31, lane 13, stream 1      
            input   wire                                        std__mgr31__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane13_strm1_data        ,
            output  wire                                        mgr31__std__lane13_strm1_data_valid  ,

            // manager 31, lane 14, stream 0      
            input   wire                                        std__mgr31__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane14_strm0_data        ,
            output  wire                                        mgr31__std__lane14_strm0_data_valid  ,

            // manager 31, lane 14, stream 1      
            input   wire                                        std__mgr31__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane14_strm1_data        ,
            output  wire                                        mgr31__std__lane14_strm1_data_valid  ,

            // manager 31, lane 15, stream 0      
            input   wire                                        std__mgr31__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane15_strm0_data        ,
            output  wire                                        mgr31__std__lane15_strm0_data_valid  ,

            // manager 31, lane 15, stream 1      
            input   wire                                        std__mgr31__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane15_strm1_data        ,
            output  wire                                        mgr31__std__lane15_strm1_data_valid  ,

            // manager 31, lane 16, stream 0      
            input   wire                                        std__mgr31__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane16_strm0_data        ,
            output  wire                                        mgr31__std__lane16_strm0_data_valid  ,

            // manager 31, lane 16, stream 1      
            input   wire                                        std__mgr31__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane16_strm1_data        ,
            output  wire                                        mgr31__std__lane16_strm1_data_valid  ,

            // manager 31, lane 17, stream 0      
            input   wire                                        std__mgr31__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane17_strm0_data        ,
            output  wire                                        mgr31__std__lane17_strm0_data_valid  ,

            // manager 31, lane 17, stream 1      
            input   wire                                        std__mgr31__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane17_strm1_data        ,
            output  wire                                        mgr31__std__lane17_strm1_data_valid  ,

            // manager 31, lane 18, stream 0      
            input   wire                                        std__mgr31__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane18_strm0_data        ,
            output  wire                                        mgr31__std__lane18_strm0_data_valid  ,

            // manager 31, lane 18, stream 1      
            input   wire                                        std__mgr31__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane18_strm1_data        ,
            output  wire                                        mgr31__std__lane18_strm1_data_valid  ,

            // manager 31, lane 19, stream 0      
            input   wire                                        std__mgr31__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane19_strm0_data        ,
            output  wire                                        mgr31__std__lane19_strm0_data_valid  ,

            // manager 31, lane 19, stream 1      
            input   wire                                        std__mgr31__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane19_strm1_data        ,
            output  wire                                        mgr31__std__lane19_strm1_data_valid  ,

            // manager 31, lane 20, stream 0      
            input   wire                                        std__mgr31__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane20_strm0_data        ,
            output  wire                                        mgr31__std__lane20_strm0_data_valid  ,

            // manager 31, lane 20, stream 1      
            input   wire                                        std__mgr31__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane20_strm1_data        ,
            output  wire                                        mgr31__std__lane20_strm1_data_valid  ,

            // manager 31, lane 21, stream 0      
            input   wire                                        std__mgr31__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane21_strm0_data        ,
            output  wire                                        mgr31__std__lane21_strm0_data_valid  ,

            // manager 31, lane 21, stream 1      
            input   wire                                        std__mgr31__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane21_strm1_data        ,
            output  wire                                        mgr31__std__lane21_strm1_data_valid  ,

            // manager 31, lane 22, stream 0      
            input   wire                                        std__mgr31__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane22_strm0_data        ,
            output  wire                                        mgr31__std__lane22_strm0_data_valid  ,

            // manager 31, lane 22, stream 1      
            input   wire                                        std__mgr31__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane22_strm1_data        ,
            output  wire                                        mgr31__std__lane22_strm1_data_valid  ,

            // manager 31, lane 23, stream 0      
            input   wire                                        std__mgr31__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane23_strm0_data        ,
            output  wire                                        mgr31__std__lane23_strm0_data_valid  ,

            // manager 31, lane 23, stream 1      
            input   wire                                        std__mgr31__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane23_strm1_data        ,
            output  wire                                        mgr31__std__lane23_strm1_data_valid  ,

            // manager 31, lane 24, stream 0      
            input   wire                                        std__mgr31__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane24_strm0_data        ,
            output  wire                                        mgr31__std__lane24_strm0_data_valid  ,

            // manager 31, lane 24, stream 1      
            input   wire                                        std__mgr31__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane24_strm1_data        ,
            output  wire                                        mgr31__std__lane24_strm1_data_valid  ,

            // manager 31, lane 25, stream 0      
            input   wire                                        std__mgr31__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane25_strm0_data        ,
            output  wire                                        mgr31__std__lane25_strm0_data_valid  ,

            // manager 31, lane 25, stream 1      
            input   wire                                        std__mgr31__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane25_strm1_data        ,
            output  wire                                        mgr31__std__lane25_strm1_data_valid  ,

            // manager 31, lane 26, stream 0      
            input   wire                                        std__mgr31__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane26_strm0_data        ,
            output  wire                                        mgr31__std__lane26_strm0_data_valid  ,

            // manager 31, lane 26, stream 1      
            input   wire                                        std__mgr31__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane26_strm1_data        ,
            output  wire                                        mgr31__std__lane26_strm1_data_valid  ,

            // manager 31, lane 27, stream 0      
            input   wire                                        std__mgr31__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane27_strm0_data        ,
            output  wire                                        mgr31__std__lane27_strm0_data_valid  ,

            // manager 31, lane 27, stream 1      
            input   wire                                        std__mgr31__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane27_strm1_data        ,
            output  wire                                        mgr31__std__lane27_strm1_data_valid  ,

            // manager 31, lane 28, stream 0      
            input   wire                                        std__mgr31__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane28_strm0_data        ,
            output  wire                                        mgr31__std__lane28_strm0_data_valid  ,

            // manager 31, lane 28, stream 1      
            input   wire                                        std__mgr31__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane28_strm1_data        ,
            output  wire                                        mgr31__std__lane28_strm1_data_valid  ,

            // manager 31, lane 29, stream 0      
            input   wire                                        std__mgr31__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane29_strm0_data        ,
            output  wire                                        mgr31__std__lane29_strm0_data_valid  ,

            // manager 31, lane 29, stream 1      
            input   wire                                        std__mgr31__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane29_strm1_data        ,
            output  wire                                        mgr31__std__lane29_strm1_data_valid  ,

            // manager 31, lane 30, stream 0      
            input   wire                                        std__mgr31__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane30_strm0_data        ,
            output  wire                                        mgr31__std__lane30_strm0_data_valid  ,

            // manager 31, lane 30, stream 1      
            input   wire                                        std__mgr31__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane30_strm1_data        ,
            output  wire                                        mgr31__std__lane30_strm1_data_valid  ,

            // manager 31, lane 31, stream 0      
            input   wire                                        std__mgr31__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane31_strm0_data        ,
            output  wire                                        mgr31__std__lane31_strm0_data_valid  ,

            // manager 31, lane 31, stream 1      
            input   wire                                        std__mgr31__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr31__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr31__std__lane31_strm1_data        ,
            output  wire                                        mgr31__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 32, lane 0, stream 0      
            input   wire                                        std__mgr32__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane0_strm0_data        ,
            output  wire                                        mgr32__std__lane0_strm0_data_valid  ,

            // manager 32, lane 0, stream 1      
            input   wire                                        std__mgr32__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane0_strm1_data        ,
            output  wire                                        mgr32__std__lane0_strm1_data_valid  ,

            // manager 32, lane 1, stream 0      
            input   wire                                        std__mgr32__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane1_strm0_data        ,
            output  wire                                        mgr32__std__lane1_strm0_data_valid  ,

            // manager 32, lane 1, stream 1      
            input   wire                                        std__mgr32__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane1_strm1_data        ,
            output  wire                                        mgr32__std__lane1_strm1_data_valid  ,

            // manager 32, lane 2, stream 0      
            input   wire                                        std__mgr32__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane2_strm0_data        ,
            output  wire                                        mgr32__std__lane2_strm0_data_valid  ,

            // manager 32, lane 2, stream 1      
            input   wire                                        std__mgr32__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane2_strm1_data        ,
            output  wire                                        mgr32__std__lane2_strm1_data_valid  ,

            // manager 32, lane 3, stream 0      
            input   wire                                        std__mgr32__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane3_strm0_data        ,
            output  wire                                        mgr32__std__lane3_strm0_data_valid  ,

            // manager 32, lane 3, stream 1      
            input   wire                                        std__mgr32__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane3_strm1_data        ,
            output  wire                                        mgr32__std__lane3_strm1_data_valid  ,

            // manager 32, lane 4, stream 0      
            input   wire                                        std__mgr32__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane4_strm0_data        ,
            output  wire                                        mgr32__std__lane4_strm0_data_valid  ,

            // manager 32, lane 4, stream 1      
            input   wire                                        std__mgr32__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane4_strm1_data        ,
            output  wire                                        mgr32__std__lane4_strm1_data_valid  ,

            // manager 32, lane 5, stream 0      
            input   wire                                        std__mgr32__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane5_strm0_data        ,
            output  wire                                        mgr32__std__lane5_strm0_data_valid  ,

            // manager 32, lane 5, stream 1      
            input   wire                                        std__mgr32__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane5_strm1_data        ,
            output  wire                                        mgr32__std__lane5_strm1_data_valid  ,

            // manager 32, lane 6, stream 0      
            input   wire                                        std__mgr32__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane6_strm0_data        ,
            output  wire                                        mgr32__std__lane6_strm0_data_valid  ,

            // manager 32, lane 6, stream 1      
            input   wire                                        std__mgr32__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane6_strm1_data        ,
            output  wire                                        mgr32__std__lane6_strm1_data_valid  ,

            // manager 32, lane 7, stream 0      
            input   wire                                        std__mgr32__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane7_strm0_data        ,
            output  wire                                        mgr32__std__lane7_strm0_data_valid  ,

            // manager 32, lane 7, stream 1      
            input   wire                                        std__mgr32__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane7_strm1_data        ,
            output  wire                                        mgr32__std__lane7_strm1_data_valid  ,

            // manager 32, lane 8, stream 0      
            input   wire                                        std__mgr32__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane8_strm0_data        ,
            output  wire                                        mgr32__std__lane8_strm0_data_valid  ,

            // manager 32, lane 8, stream 1      
            input   wire                                        std__mgr32__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane8_strm1_data        ,
            output  wire                                        mgr32__std__lane8_strm1_data_valid  ,

            // manager 32, lane 9, stream 0      
            input   wire                                        std__mgr32__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane9_strm0_data        ,
            output  wire                                        mgr32__std__lane9_strm0_data_valid  ,

            // manager 32, lane 9, stream 1      
            input   wire                                        std__mgr32__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane9_strm1_data        ,
            output  wire                                        mgr32__std__lane9_strm1_data_valid  ,

            // manager 32, lane 10, stream 0      
            input   wire                                        std__mgr32__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane10_strm0_data        ,
            output  wire                                        mgr32__std__lane10_strm0_data_valid  ,

            // manager 32, lane 10, stream 1      
            input   wire                                        std__mgr32__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane10_strm1_data        ,
            output  wire                                        mgr32__std__lane10_strm1_data_valid  ,

            // manager 32, lane 11, stream 0      
            input   wire                                        std__mgr32__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane11_strm0_data        ,
            output  wire                                        mgr32__std__lane11_strm0_data_valid  ,

            // manager 32, lane 11, stream 1      
            input   wire                                        std__mgr32__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane11_strm1_data        ,
            output  wire                                        mgr32__std__lane11_strm1_data_valid  ,

            // manager 32, lane 12, stream 0      
            input   wire                                        std__mgr32__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane12_strm0_data        ,
            output  wire                                        mgr32__std__lane12_strm0_data_valid  ,

            // manager 32, lane 12, stream 1      
            input   wire                                        std__mgr32__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane12_strm1_data        ,
            output  wire                                        mgr32__std__lane12_strm1_data_valid  ,

            // manager 32, lane 13, stream 0      
            input   wire                                        std__mgr32__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane13_strm0_data        ,
            output  wire                                        mgr32__std__lane13_strm0_data_valid  ,

            // manager 32, lane 13, stream 1      
            input   wire                                        std__mgr32__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane13_strm1_data        ,
            output  wire                                        mgr32__std__lane13_strm1_data_valid  ,

            // manager 32, lane 14, stream 0      
            input   wire                                        std__mgr32__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane14_strm0_data        ,
            output  wire                                        mgr32__std__lane14_strm0_data_valid  ,

            // manager 32, lane 14, stream 1      
            input   wire                                        std__mgr32__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane14_strm1_data        ,
            output  wire                                        mgr32__std__lane14_strm1_data_valid  ,

            // manager 32, lane 15, stream 0      
            input   wire                                        std__mgr32__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane15_strm0_data        ,
            output  wire                                        mgr32__std__lane15_strm0_data_valid  ,

            // manager 32, lane 15, stream 1      
            input   wire                                        std__mgr32__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane15_strm1_data        ,
            output  wire                                        mgr32__std__lane15_strm1_data_valid  ,

            // manager 32, lane 16, stream 0      
            input   wire                                        std__mgr32__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane16_strm0_data        ,
            output  wire                                        mgr32__std__lane16_strm0_data_valid  ,

            // manager 32, lane 16, stream 1      
            input   wire                                        std__mgr32__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane16_strm1_data        ,
            output  wire                                        mgr32__std__lane16_strm1_data_valid  ,

            // manager 32, lane 17, stream 0      
            input   wire                                        std__mgr32__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane17_strm0_data        ,
            output  wire                                        mgr32__std__lane17_strm0_data_valid  ,

            // manager 32, lane 17, stream 1      
            input   wire                                        std__mgr32__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane17_strm1_data        ,
            output  wire                                        mgr32__std__lane17_strm1_data_valid  ,

            // manager 32, lane 18, stream 0      
            input   wire                                        std__mgr32__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane18_strm0_data        ,
            output  wire                                        mgr32__std__lane18_strm0_data_valid  ,

            // manager 32, lane 18, stream 1      
            input   wire                                        std__mgr32__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane18_strm1_data        ,
            output  wire                                        mgr32__std__lane18_strm1_data_valid  ,

            // manager 32, lane 19, stream 0      
            input   wire                                        std__mgr32__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane19_strm0_data        ,
            output  wire                                        mgr32__std__lane19_strm0_data_valid  ,

            // manager 32, lane 19, stream 1      
            input   wire                                        std__mgr32__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane19_strm1_data        ,
            output  wire                                        mgr32__std__lane19_strm1_data_valid  ,

            // manager 32, lane 20, stream 0      
            input   wire                                        std__mgr32__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane20_strm0_data        ,
            output  wire                                        mgr32__std__lane20_strm0_data_valid  ,

            // manager 32, lane 20, stream 1      
            input   wire                                        std__mgr32__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane20_strm1_data        ,
            output  wire                                        mgr32__std__lane20_strm1_data_valid  ,

            // manager 32, lane 21, stream 0      
            input   wire                                        std__mgr32__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane21_strm0_data        ,
            output  wire                                        mgr32__std__lane21_strm0_data_valid  ,

            // manager 32, lane 21, stream 1      
            input   wire                                        std__mgr32__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane21_strm1_data        ,
            output  wire                                        mgr32__std__lane21_strm1_data_valid  ,

            // manager 32, lane 22, stream 0      
            input   wire                                        std__mgr32__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane22_strm0_data        ,
            output  wire                                        mgr32__std__lane22_strm0_data_valid  ,

            // manager 32, lane 22, stream 1      
            input   wire                                        std__mgr32__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane22_strm1_data        ,
            output  wire                                        mgr32__std__lane22_strm1_data_valid  ,

            // manager 32, lane 23, stream 0      
            input   wire                                        std__mgr32__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane23_strm0_data        ,
            output  wire                                        mgr32__std__lane23_strm0_data_valid  ,

            // manager 32, lane 23, stream 1      
            input   wire                                        std__mgr32__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane23_strm1_data        ,
            output  wire                                        mgr32__std__lane23_strm1_data_valid  ,

            // manager 32, lane 24, stream 0      
            input   wire                                        std__mgr32__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane24_strm0_data        ,
            output  wire                                        mgr32__std__lane24_strm0_data_valid  ,

            // manager 32, lane 24, stream 1      
            input   wire                                        std__mgr32__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane24_strm1_data        ,
            output  wire                                        mgr32__std__lane24_strm1_data_valid  ,

            // manager 32, lane 25, stream 0      
            input   wire                                        std__mgr32__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane25_strm0_data        ,
            output  wire                                        mgr32__std__lane25_strm0_data_valid  ,

            // manager 32, lane 25, stream 1      
            input   wire                                        std__mgr32__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane25_strm1_data        ,
            output  wire                                        mgr32__std__lane25_strm1_data_valid  ,

            // manager 32, lane 26, stream 0      
            input   wire                                        std__mgr32__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane26_strm0_data        ,
            output  wire                                        mgr32__std__lane26_strm0_data_valid  ,

            // manager 32, lane 26, stream 1      
            input   wire                                        std__mgr32__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane26_strm1_data        ,
            output  wire                                        mgr32__std__lane26_strm1_data_valid  ,

            // manager 32, lane 27, stream 0      
            input   wire                                        std__mgr32__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane27_strm0_data        ,
            output  wire                                        mgr32__std__lane27_strm0_data_valid  ,

            // manager 32, lane 27, stream 1      
            input   wire                                        std__mgr32__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane27_strm1_data        ,
            output  wire                                        mgr32__std__lane27_strm1_data_valid  ,

            // manager 32, lane 28, stream 0      
            input   wire                                        std__mgr32__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane28_strm0_data        ,
            output  wire                                        mgr32__std__lane28_strm0_data_valid  ,

            // manager 32, lane 28, stream 1      
            input   wire                                        std__mgr32__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane28_strm1_data        ,
            output  wire                                        mgr32__std__lane28_strm1_data_valid  ,

            // manager 32, lane 29, stream 0      
            input   wire                                        std__mgr32__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane29_strm0_data        ,
            output  wire                                        mgr32__std__lane29_strm0_data_valid  ,

            // manager 32, lane 29, stream 1      
            input   wire                                        std__mgr32__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane29_strm1_data        ,
            output  wire                                        mgr32__std__lane29_strm1_data_valid  ,

            // manager 32, lane 30, stream 0      
            input   wire                                        std__mgr32__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane30_strm0_data        ,
            output  wire                                        mgr32__std__lane30_strm0_data_valid  ,

            // manager 32, lane 30, stream 1      
            input   wire                                        std__mgr32__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane30_strm1_data        ,
            output  wire                                        mgr32__std__lane30_strm1_data_valid  ,

            // manager 32, lane 31, stream 0      
            input   wire                                        std__mgr32__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane31_strm0_data        ,
            output  wire                                        mgr32__std__lane31_strm0_data_valid  ,

            // manager 32, lane 31, stream 1      
            input   wire                                        std__mgr32__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr32__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr32__std__lane31_strm1_data        ,
            output  wire                                        mgr32__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 33, lane 0, stream 0      
            input   wire                                        std__mgr33__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane0_strm0_data        ,
            output  wire                                        mgr33__std__lane0_strm0_data_valid  ,

            // manager 33, lane 0, stream 1      
            input   wire                                        std__mgr33__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane0_strm1_data        ,
            output  wire                                        mgr33__std__lane0_strm1_data_valid  ,

            // manager 33, lane 1, stream 0      
            input   wire                                        std__mgr33__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane1_strm0_data        ,
            output  wire                                        mgr33__std__lane1_strm0_data_valid  ,

            // manager 33, lane 1, stream 1      
            input   wire                                        std__mgr33__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane1_strm1_data        ,
            output  wire                                        mgr33__std__lane1_strm1_data_valid  ,

            // manager 33, lane 2, stream 0      
            input   wire                                        std__mgr33__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane2_strm0_data        ,
            output  wire                                        mgr33__std__lane2_strm0_data_valid  ,

            // manager 33, lane 2, stream 1      
            input   wire                                        std__mgr33__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane2_strm1_data        ,
            output  wire                                        mgr33__std__lane2_strm1_data_valid  ,

            // manager 33, lane 3, stream 0      
            input   wire                                        std__mgr33__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane3_strm0_data        ,
            output  wire                                        mgr33__std__lane3_strm0_data_valid  ,

            // manager 33, lane 3, stream 1      
            input   wire                                        std__mgr33__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane3_strm1_data        ,
            output  wire                                        mgr33__std__lane3_strm1_data_valid  ,

            // manager 33, lane 4, stream 0      
            input   wire                                        std__mgr33__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane4_strm0_data        ,
            output  wire                                        mgr33__std__lane4_strm0_data_valid  ,

            // manager 33, lane 4, stream 1      
            input   wire                                        std__mgr33__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane4_strm1_data        ,
            output  wire                                        mgr33__std__lane4_strm1_data_valid  ,

            // manager 33, lane 5, stream 0      
            input   wire                                        std__mgr33__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane5_strm0_data        ,
            output  wire                                        mgr33__std__lane5_strm0_data_valid  ,

            // manager 33, lane 5, stream 1      
            input   wire                                        std__mgr33__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane5_strm1_data        ,
            output  wire                                        mgr33__std__lane5_strm1_data_valid  ,

            // manager 33, lane 6, stream 0      
            input   wire                                        std__mgr33__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane6_strm0_data        ,
            output  wire                                        mgr33__std__lane6_strm0_data_valid  ,

            // manager 33, lane 6, stream 1      
            input   wire                                        std__mgr33__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane6_strm1_data        ,
            output  wire                                        mgr33__std__lane6_strm1_data_valid  ,

            // manager 33, lane 7, stream 0      
            input   wire                                        std__mgr33__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane7_strm0_data        ,
            output  wire                                        mgr33__std__lane7_strm0_data_valid  ,

            // manager 33, lane 7, stream 1      
            input   wire                                        std__mgr33__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane7_strm1_data        ,
            output  wire                                        mgr33__std__lane7_strm1_data_valid  ,

            // manager 33, lane 8, stream 0      
            input   wire                                        std__mgr33__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane8_strm0_data        ,
            output  wire                                        mgr33__std__lane8_strm0_data_valid  ,

            // manager 33, lane 8, stream 1      
            input   wire                                        std__mgr33__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane8_strm1_data        ,
            output  wire                                        mgr33__std__lane8_strm1_data_valid  ,

            // manager 33, lane 9, stream 0      
            input   wire                                        std__mgr33__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane9_strm0_data        ,
            output  wire                                        mgr33__std__lane9_strm0_data_valid  ,

            // manager 33, lane 9, stream 1      
            input   wire                                        std__mgr33__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane9_strm1_data        ,
            output  wire                                        mgr33__std__lane9_strm1_data_valid  ,

            // manager 33, lane 10, stream 0      
            input   wire                                        std__mgr33__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane10_strm0_data        ,
            output  wire                                        mgr33__std__lane10_strm0_data_valid  ,

            // manager 33, lane 10, stream 1      
            input   wire                                        std__mgr33__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane10_strm1_data        ,
            output  wire                                        mgr33__std__lane10_strm1_data_valid  ,

            // manager 33, lane 11, stream 0      
            input   wire                                        std__mgr33__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane11_strm0_data        ,
            output  wire                                        mgr33__std__lane11_strm0_data_valid  ,

            // manager 33, lane 11, stream 1      
            input   wire                                        std__mgr33__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane11_strm1_data        ,
            output  wire                                        mgr33__std__lane11_strm1_data_valid  ,

            // manager 33, lane 12, stream 0      
            input   wire                                        std__mgr33__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane12_strm0_data        ,
            output  wire                                        mgr33__std__lane12_strm0_data_valid  ,

            // manager 33, lane 12, stream 1      
            input   wire                                        std__mgr33__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane12_strm1_data        ,
            output  wire                                        mgr33__std__lane12_strm1_data_valid  ,

            // manager 33, lane 13, stream 0      
            input   wire                                        std__mgr33__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane13_strm0_data        ,
            output  wire                                        mgr33__std__lane13_strm0_data_valid  ,

            // manager 33, lane 13, stream 1      
            input   wire                                        std__mgr33__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane13_strm1_data        ,
            output  wire                                        mgr33__std__lane13_strm1_data_valid  ,

            // manager 33, lane 14, stream 0      
            input   wire                                        std__mgr33__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane14_strm0_data        ,
            output  wire                                        mgr33__std__lane14_strm0_data_valid  ,

            // manager 33, lane 14, stream 1      
            input   wire                                        std__mgr33__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane14_strm1_data        ,
            output  wire                                        mgr33__std__lane14_strm1_data_valid  ,

            // manager 33, lane 15, stream 0      
            input   wire                                        std__mgr33__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane15_strm0_data        ,
            output  wire                                        mgr33__std__lane15_strm0_data_valid  ,

            // manager 33, lane 15, stream 1      
            input   wire                                        std__mgr33__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane15_strm1_data        ,
            output  wire                                        mgr33__std__lane15_strm1_data_valid  ,

            // manager 33, lane 16, stream 0      
            input   wire                                        std__mgr33__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane16_strm0_data        ,
            output  wire                                        mgr33__std__lane16_strm0_data_valid  ,

            // manager 33, lane 16, stream 1      
            input   wire                                        std__mgr33__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane16_strm1_data        ,
            output  wire                                        mgr33__std__lane16_strm1_data_valid  ,

            // manager 33, lane 17, stream 0      
            input   wire                                        std__mgr33__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane17_strm0_data        ,
            output  wire                                        mgr33__std__lane17_strm0_data_valid  ,

            // manager 33, lane 17, stream 1      
            input   wire                                        std__mgr33__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane17_strm1_data        ,
            output  wire                                        mgr33__std__lane17_strm1_data_valid  ,

            // manager 33, lane 18, stream 0      
            input   wire                                        std__mgr33__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane18_strm0_data        ,
            output  wire                                        mgr33__std__lane18_strm0_data_valid  ,

            // manager 33, lane 18, stream 1      
            input   wire                                        std__mgr33__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane18_strm1_data        ,
            output  wire                                        mgr33__std__lane18_strm1_data_valid  ,

            // manager 33, lane 19, stream 0      
            input   wire                                        std__mgr33__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane19_strm0_data        ,
            output  wire                                        mgr33__std__lane19_strm0_data_valid  ,

            // manager 33, lane 19, stream 1      
            input   wire                                        std__mgr33__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane19_strm1_data        ,
            output  wire                                        mgr33__std__lane19_strm1_data_valid  ,

            // manager 33, lane 20, stream 0      
            input   wire                                        std__mgr33__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane20_strm0_data        ,
            output  wire                                        mgr33__std__lane20_strm0_data_valid  ,

            // manager 33, lane 20, stream 1      
            input   wire                                        std__mgr33__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane20_strm1_data        ,
            output  wire                                        mgr33__std__lane20_strm1_data_valid  ,

            // manager 33, lane 21, stream 0      
            input   wire                                        std__mgr33__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane21_strm0_data        ,
            output  wire                                        mgr33__std__lane21_strm0_data_valid  ,

            // manager 33, lane 21, stream 1      
            input   wire                                        std__mgr33__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane21_strm1_data        ,
            output  wire                                        mgr33__std__lane21_strm1_data_valid  ,

            // manager 33, lane 22, stream 0      
            input   wire                                        std__mgr33__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane22_strm0_data        ,
            output  wire                                        mgr33__std__lane22_strm0_data_valid  ,

            // manager 33, lane 22, stream 1      
            input   wire                                        std__mgr33__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane22_strm1_data        ,
            output  wire                                        mgr33__std__lane22_strm1_data_valid  ,

            // manager 33, lane 23, stream 0      
            input   wire                                        std__mgr33__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane23_strm0_data        ,
            output  wire                                        mgr33__std__lane23_strm0_data_valid  ,

            // manager 33, lane 23, stream 1      
            input   wire                                        std__mgr33__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane23_strm1_data        ,
            output  wire                                        mgr33__std__lane23_strm1_data_valid  ,

            // manager 33, lane 24, stream 0      
            input   wire                                        std__mgr33__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane24_strm0_data        ,
            output  wire                                        mgr33__std__lane24_strm0_data_valid  ,

            // manager 33, lane 24, stream 1      
            input   wire                                        std__mgr33__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane24_strm1_data        ,
            output  wire                                        mgr33__std__lane24_strm1_data_valid  ,

            // manager 33, lane 25, stream 0      
            input   wire                                        std__mgr33__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane25_strm0_data        ,
            output  wire                                        mgr33__std__lane25_strm0_data_valid  ,

            // manager 33, lane 25, stream 1      
            input   wire                                        std__mgr33__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane25_strm1_data        ,
            output  wire                                        mgr33__std__lane25_strm1_data_valid  ,

            // manager 33, lane 26, stream 0      
            input   wire                                        std__mgr33__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane26_strm0_data        ,
            output  wire                                        mgr33__std__lane26_strm0_data_valid  ,

            // manager 33, lane 26, stream 1      
            input   wire                                        std__mgr33__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane26_strm1_data        ,
            output  wire                                        mgr33__std__lane26_strm1_data_valid  ,

            // manager 33, lane 27, stream 0      
            input   wire                                        std__mgr33__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane27_strm0_data        ,
            output  wire                                        mgr33__std__lane27_strm0_data_valid  ,

            // manager 33, lane 27, stream 1      
            input   wire                                        std__mgr33__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane27_strm1_data        ,
            output  wire                                        mgr33__std__lane27_strm1_data_valid  ,

            // manager 33, lane 28, stream 0      
            input   wire                                        std__mgr33__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane28_strm0_data        ,
            output  wire                                        mgr33__std__lane28_strm0_data_valid  ,

            // manager 33, lane 28, stream 1      
            input   wire                                        std__mgr33__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane28_strm1_data        ,
            output  wire                                        mgr33__std__lane28_strm1_data_valid  ,

            // manager 33, lane 29, stream 0      
            input   wire                                        std__mgr33__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane29_strm0_data        ,
            output  wire                                        mgr33__std__lane29_strm0_data_valid  ,

            // manager 33, lane 29, stream 1      
            input   wire                                        std__mgr33__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane29_strm1_data        ,
            output  wire                                        mgr33__std__lane29_strm1_data_valid  ,

            // manager 33, lane 30, stream 0      
            input   wire                                        std__mgr33__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane30_strm0_data        ,
            output  wire                                        mgr33__std__lane30_strm0_data_valid  ,

            // manager 33, lane 30, stream 1      
            input   wire                                        std__mgr33__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane30_strm1_data        ,
            output  wire                                        mgr33__std__lane30_strm1_data_valid  ,

            // manager 33, lane 31, stream 0      
            input   wire                                        std__mgr33__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane31_strm0_data        ,
            output  wire                                        mgr33__std__lane31_strm0_data_valid  ,

            // manager 33, lane 31, stream 1      
            input   wire                                        std__mgr33__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr33__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr33__std__lane31_strm1_data        ,
            output  wire                                        mgr33__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 34, lane 0, stream 0      
            input   wire                                        std__mgr34__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane0_strm0_data        ,
            output  wire                                        mgr34__std__lane0_strm0_data_valid  ,

            // manager 34, lane 0, stream 1      
            input   wire                                        std__mgr34__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane0_strm1_data        ,
            output  wire                                        mgr34__std__lane0_strm1_data_valid  ,

            // manager 34, lane 1, stream 0      
            input   wire                                        std__mgr34__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane1_strm0_data        ,
            output  wire                                        mgr34__std__lane1_strm0_data_valid  ,

            // manager 34, lane 1, stream 1      
            input   wire                                        std__mgr34__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane1_strm1_data        ,
            output  wire                                        mgr34__std__lane1_strm1_data_valid  ,

            // manager 34, lane 2, stream 0      
            input   wire                                        std__mgr34__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane2_strm0_data        ,
            output  wire                                        mgr34__std__lane2_strm0_data_valid  ,

            // manager 34, lane 2, stream 1      
            input   wire                                        std__mgr34__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane2_strm1_data        ,
            output  wire                                        mgr34__std__lane2_strm1_data_valid  ,

            // manager 34, lane 3, stream 0      
            input   wire                                        std__mgr34__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane3_strm0_data        ,
            output  wire                                        mgr34__std__lane3_strm0_data_valid  ,

            // manager 34, lane 3, stream 1      
            input   wire                                        std__mgr34__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane3_strm1_data        ,
            output  wire                                        mgr34__std__lane3_strm1_data_valid  ,

            // manager 34, lane 4, stream 0      
            input   wire                                        std__mgr34__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane4_strm0_data        ,
            output  wire                                        mgr34__std__lane4_strm0_data_valid  ,

            // manager 34, lane 4, stream 1      
            input   wire                                        std__mgr34__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane4_strm1_data        ,
            output  wire                                        mgr34__std__lane4_strm1_data_valid  ,

            // manager 34, lane 5, stream 0      
            input   wire                                        std__mgr34__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane5_strm0_data        ,
            output  wire                                        mgr34__std__lane5_strm0_data_valid  ,

            // manager 34, lane 5, stream 1      
            input   wire                                        std__mgr34__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane5_strm1_data        ,
            output  wire                                        mgr34__std__lane5_strm1_data_valid  ,

            // manager 34, lane 6, stream 0      
            input   wire                                        std__mgr34__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane6_strm0_data        ,
            output  wire                                        mgr34__std__lane6_strm0_data_valid  ,

            // manager 34, lane 6, stream 1      
            input   wire                                        std__mgr34__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane6_strm1_data        ,
            output  wire                                        mgr34__std__lane6_strm1_data_valid  ,

            // manager 34, lane 7, stream 0      
            input   wire                                        std__mgr34__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane7_strm0_data        ,
            output  wire                                        mgr34__std__lane7_strm0_data_valid  ,

            // manager 34, lane 7, stream 1      
            input   wire                                        std__mgr34__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane7_strm1_data        ,
            output  wire                                        mgr34__std__lane7_strm1_data_valid  ,

            // manager 34, lane 8, stream 0      
            input   wire                                        std__mgr34__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane8_strm0_data        ,
            output  wire                                        mgr34__std__lane8_strm0_data_valid  ,

            // manager 34, lane 8, stream 1      
            input   wire                                        std__mgr34__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane8_strm1_data        ,
            output  wire                                        mgr34__std__lane8_strm1_data_valid  ,

            // manager 34, lane 9, stream 0      
            input   wire                                        std__mgr34__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane9_strm0_data        ,
            output  wire                                        mgr34__std__lane9_strm0_data_valid  ,

            // manager 34, lane 9, stream 1      
            input   wire                                        std__mgr34__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane9_strm1_data        ,
            output  wire                                        mgr34__std__lane9_strm1_data_valid  ,

            // manager 34, lane 10, stream 0      
            input   wire                                        std__mgr34__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane10_strm0_data        ,
            output  wire                                        mgr34__std__lane10_strm0_data_valid  ,

            // manager 34, lane 10, stream 1      
            input   wire                                        std__mgr34__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane10_strm1_data        ,
            output  wire                                        mgr34__std__lane10_strm1_data_valid  ,

            // manager 34, lane 11, stream 0      
            input   wire                                        std__mgr34__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane11_strm0_data        ,
            output  wire                                        mgr34__std__lane11_strm0_data_valid  ,

            // manager 34, lane 11, stream 1      
            input   wire                                        std__mgr34__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane11_strm1_data        ,
            output  wire                                        mgr34__std__lane11_strm1_data_valid  ,

            // manager 34, lane 12, stream 0      
            input   wire                                        std__mgr34__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane12_strm0_data        ,
            output  wire                                        mgr34__std__lane12_strm0_data_valid  ,

            // manager 34, lane 12, stream 1      
            input   wire                                        std__mgr34__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane12_strm1_data        ,
            output  wire                                        mgr34__std__lane12_strm1_data_valid  ,

            // manager 34, lane 13, stream 0      
            input   wire                                        std__mgr34__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane13_strm0_data        ,
            output  wire                                        mgr34__std__lane13_strm0_data_valid  ,

            // manager 34, lane 13, stream 1      
            input   wire                                        std__mgr34__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane13_strm1_data        ,
            output  wire                                        mgr34__std__lane13_strm1_data_valid  ,

            // manager 34, lane 14, stream 0      
            input   wire                                        std__mgr34__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane14_strm0_data        ,
            output  wire                                        mgr34__std__lane14_strm0_data_valid  ,

            // manager 34, lane 14, stream 1      
            input   wire                                        std__mgr34__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane14_strm1_data        ,
            output  wire                                        mgr34__std__lane14_strm1_data_valid  ,

            // manager 34, lane 15, stream 0      
            input   wire                                        std__mgr34__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane15_strm0_data        ,
            output  wire                                        mgr34__std__lane15_strm0_data_valid  ,

            // manager 34, lane 15, stream 1      
            input   wire                                        std__mgr34__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane15_strm1_data        ,
            output  wire                                        mgr34__std__lane15_strm1_data_valid  ,

            // manager 34, lane 16, stream 0      
            input   wire                                        std__mgr34__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane16_strm0_data        ,
            output  wire                                        mgr34__std__lane16_strm0_data_valid  ,

            // manager 34, lane 16, stream 1      
            input   wire                                        std__mgr34__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane16_strm1_data        ,
            output  wire                                        mgr34__std__lane16_strm1_data_valid  ,

            // manager 34, lane 17, stream 0      
            input   wire                                        std__mgr34__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane17_strm0_data        ,
            output  wire                                        mgr34__std__lane17_strm0_data_valid  ,

            // manager 34, lane 17, stream 1      
            input   wire                                        std__mgr34__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane17_strm1_data        ,
            output  wire                                        mgr34__std__lane17_strm1_data_valid  ,

            // manager 34, lane 18, stream 0      
            input   wire                                        std__mgr34__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane18_strm0_data        ,
            output  wire                                        mgr34__std__lane18_strm0_data_valid  ,

            // manager 34, lane 18, stream 1      
            input   wire                                        std__mgr34__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane18_strm1_data        ,
            output  wire                                        mgr34__std__lane18_strm1_data_valid  ,

            // manager 34, lane 19, stream 0      
            input   wire                                        std__mgr34__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane19_strm0_data        ,
            output  wire                                        mgr34__std__lane19_strm0_data_valid  ,

            // manager 34, lane 19, stream 1      
            input   wire                                        std__mgr34__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane19_strm1_data        ,
            output  wire                                        mgr34__std__lane19_strm1_data_valid  ,

            // manager 34, lane 20, stream 0      
            input   wire                                        std__mgr34__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane20_strm0_data        ,
            output  wire                                        mgr34__std__lane20_strm0_data_valid  ,

            // manager 34, lane 20, stream 1      
            input   wire                                        std__mgr34__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane20_strm1_data        ,
            output  wire                                        mgr34__std__lane20_strm1_data_valid  ,

            // manager 34, lane 21, stream 0      
            input   wire                                        std__mgr34__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane21_strm0_data        ,
            output  wire                                        mgr34__std__lane21_strm0_data_valid  ,

            // manager 34, lane 21, stream 1      
            input   wire                                        std__mgr34__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane21_strm1_data        ,
            output  wire                                        mgr34__std__lane21_strm1_data_valid  ,

            // manager 34, lane 22, stream 0      
            input   wire                                        std__mgr34__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane22_strm0_data        ,
            output  wire                                        mgr34__std__lane22_strm0_data_valid  ,

            // manager 34, lane 22, stream 1      
            input   wire                                        std__mgr34__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane22_strm1_data        ,
            output  wire                                        mgr34__std__lane22_strm1_data_valid  ,

            // manager 34, lane 23, stream 0      
            input   wire                                        std__mgr34__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane23_strm0_data        ,
            output  wire                                        mgr34__std__lane23_strm0_data_valid  ,

            // manager 34, lane 23, stream 1      
            input   wire                                        std__mgr34__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane23_strm1_data        ,
            output  wire                                        mgr34__std__lane23_strm1_data_valid  ,

            // manager 34, lane 24, stream 0      
            input   wire                                        std__mgr34__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane24_strm0_data        ,
            output  wire                                        mgr34__std__lane24_strm0_data_valid  ,

            // manager 34, lane 24, stream 1      
            input   wire                                        std__mgr34__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane24_strm1_data        ,
            output  wire                                        mgr34__std__lane24_strm1_data_valid  ,

            // manager 34, lane 25, stream 0      
            input   wire                                        std__mgr34__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane25_strm0_data        ,
            output  wire                                        mgr34__std__lane25_strm0_data_valid  ,

            // manager 34, lane 25, stream 1      
            input   wire                                        std__mgr34__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane25_strm1_data        ,
            output  wire                                        mgr34__std__lane25_strm1_data_valid  ,

            // manager 34, lane 26, stream 0      
            input   wire                                        std__mgr34__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane26_strm0_data        ,
            output  wire                                        mgr34__std__lane26_strm0_data_valid  ,

            // manager 34, lane 26, stream 1      
            input   wire                                        std__mgr34__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane26_strm1_data        ,
            output  wire                                        mgr34__std__lane26_strm1_data_valid  ,

            // manager 34, lane 27, stream 0      
            input   wire                                        std__mgr34__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane27_strm0_data        ,
            output  wire                                        mgr34__std__lane27_strm0_data_valid  ,

            // manager 34, lane 27, stream 1      
            input   wire                                        std__mgr34__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane27_strm1_data        ,
            output  wire                                        mgr34__std__lane27_strm1_data_valid  ,

            // manager 34, lane 28, stream 0      
            input   wire                                        std__mgr34__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane28_strm0_data        ,
            output  wire                                        mgr34__std__lane28_strm0_data_valid  ,

            // manager 34, lane 28, stream 1      
            input   wire                                        std__mgr34__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane28_strm1_data        ,
            output  wire                                        mgr34__std__lane28_strm1_data_valid  ,

            // manager 34, lane 29, stream 0      
            input   wire                                        std__mgr34__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane29_strm0_data        ,
            output  wire                                        mgr34__std__lane29_strm0_data_valid  ,

            // manager 34, lane 29, stream 1      
            input   wire                                        std__mgr34__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane29_strm1_data        ,
            output  wire                                        mgr34__std__lane29_strm1_data_valid  ,

            // manager 34, lane 30, stream 0      
            input   wire                                        std__mgr34__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane30_strm0_data        ,
            output  wire                                        mgr34__std__lane30_strm0_data_valid  ,

            // manager 34, lane 30, stream 1      
            input   wire                                        std__mgr34__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane30_strm1_data        ,
            output  wire                                        mgr34__std__lane30_strm1_data_valid  ,

            // manager 34, lane 31, stream 0      
            input   wire                                        std__mgr34__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane31_strm0_data        ,
            output  wire                                        mgr34__std__lane31_strm0_data_valid  ,

            // manager 34, lane 31, stream 1      
            input   wire                                        std__mgr34__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr34__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr34__std__lane31_strm1_data        ,
            output  wire                                        mgr34__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 35, lane 0, stream 0      
            input   wire                                        std__mgr35__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane0_strm0_data        ,
            output  wire                                        mgr35__std__lane0_strm0_data_valid  ,

            // manager 35, lane 0, stream 1      
            input   wire                                        std__mgr35__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane0_strm1_data        ,
            output  wire                                        mgr35__std__lane0_strm1_data_valid  ,

            // manager 35, lane 1, stream 0      
            input   wire                                        std__mgr35__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane1_strm0_data        ,
            output  wire                                        mgr35__std__lane1_strm0_data_valid  ,

            // manager 35, lane 1, stream 1      
            input   wire                                        std__mgr35__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane1_strm1_data        ,
            output  wire                                        mgr35__std__lane1_strm1_data_valid  ,

            // manager 35, lane 2, stream 0      
            input   wire                                        std__mgr35__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane2_strm0_data        ,
            output  wire                                        mgr35__std__lane2_strm0_data_valid  ,

            // manager 35, lane 2, stream 1      
            input   wire                                        std__mgr35__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane2_strm1_data        ,
            output  wire                                        mgr35__std__lane2_strm1_data_valid  ,

            // manager 35, lane 3, stream 0      
            input   wire                                        std__mgr35__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane3_strm0_data        ,
            output  wire                                        mgr35__std__lane3_strm0_data_valid  ,

            // manager 35, lane 3, stream 1      
            input   wire                                        std__mgr35__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane3_strm1_data        ,
            output  wire                                        mgr35__std__lane3_strm1_data_valid  ,

            // manager 35, lane 4, stream 0      
            input   wire                                        std__mgr35__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane4_strm0_data        ,
            output  wire                                        mgr35__std__lane4_strm0_data_valid  ,

            // manager 35, lane 4, stream 1      
            input   wire                                        std__mgr35__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane4_strm1_data        ,
            output  wire                                        mgr35__std__lane4_strm1_data_valid  ,

            // manager 35, lane 5, stream 0      
            input   wire                                        std__mgr35__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane5_strm0_data        ,
            output  wire                                        mgr35__std__lane5_strm0_data_valid  ,

            // manager 35, lane 5, stream 1      
            input   wire                                        std__mgr35__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane5_strm1_data        ,
            output  wire                                        mgr35__std__lane5_strm1_data_valid  ,

            // manager 35, lane 6, stream 0      
            input   wire                                        std__mgr35__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane6_strm0_data        ,
            output  wire                                        mgr35__std__lane6_strm0_data_valid  ,

            // manager 35, lane 6, stream 1      
            input   wire                                        std__mgr35__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane6_strm1_data        ,
            output  wire                                        mgr35__std__lane6_strm1_data_valid  ,

            // manager 35, lane 7, stream 0      
            input   wire                                        std__mgr35__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane7_strm0_data        ,
            output  wire                                        mgr35__std__lane7_strm0_data_valid  ,

            // manager 35, lane 7, stream 1      
            input   wire                                        std__mgr35__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane7_strm1_data        ,
            output  wire                                        mgr35__std__lane7_strm1_data_valid  ,

            // manager 35, lane 8, stream 0      
            input   wire                                        std__mgr35__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane8_strm0_data        ,
            output  wire                                        mgr35__std__lane8_strm0_data_valid  ,

            // manager 35, lane 8, stream 1      
            input   wire                                        std__mgr35__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane8_strm1_data        ,
            output  wire                                        mgr35__std__lane8_strm1_data_valid  ,

            // manager 35, lane 9, stream 0      
            input   wire                                        std__mgr35__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane9_strm0_data        ,
            output  wire                                        mgr35__std__lane9_strm0_data_valid  ,

            // manager 35, lane 9, stream 1      
            input   wire                                        std__mgr35__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane9_strm1_data        ,
            output  wire                                        mgr35__std__lane9_strm1_data_valid  ,

            // manager 35, lane 10, stream 0      
            input   wire                                        std__mgr35__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane10_strm0_data        ,
            output  wire                                        mgr35__std__lane10_strm0_data_valid  ,

            // manager 35, lane 10, stream 1      
            input   wire                                        std__mgr35__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane10_strm1_data        ,
            output  wire                                        mgr35__std__lane10_strm1_data_valid  ,

            // manager 35, lane 11, stream 0      
            input   wire                                        std__mgr35__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane11_strm0_data        ,
            output  wire                                        mgr35__std__lane11_strm0_data_valid  ,

            // manager 35, lane 11, stream 1      
            input   wire                                        std__mgr35__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane11_strm1_data        ,
            output  wire                                        mgr35__std__lane11_strm1_data_valid  ,

            // manager 35, lane 12, stream 0      
            input   wire                                        std__mgr35__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane12_strm0_data        ,
            output  wire                                        mgr35__std__lane12_strm0_data_valid  ,

            // manager 35, lane 12, stream 1      
            input   wire                                        std__mgr35__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane12_strm1_data        ,
            output  wire                                        mgr35__std__lane12_strm1_data_valid  ,

            // manager 35, lane 13, stream 0      
            input   wire                                        std__mgr35__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane13_strm0_data        ,
            output  wire                                        mgr35__std__lane13_strm0_data_valid  ,

            // manager 35, lane 13, stream 1      
            input   wire                                        std__mgr35__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane13_strm1_data        ,
            output  wire                                        mgr35__std__lane13_strm1_data_valid  ,

            // manager 35, lane 14, stream 0      
            input   wire                                        std__mgr35__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane14_strm0_data        ,
            output  wire                                        mgr35__std__lane14_strm0_data_valid  ,

            // manager 35, lane 14, stream 1      
            input   wire                                        std__mgr35__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane14_strm1_data        ,
            output  wire                                        mgr35__std__lane14_strm1_data_valid  ,

            // manager 35, lane 15, stream 0      
            input   wire                                        std__mgr35__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane15_strm0_data        ,
            output  wire                                        mgr35__std__lane15_strm0_data_valid  ,

            // manager 35, lane 15, stream 1      
            input   wire                                        std__mgr35__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane15_strm1_data        ,
            output  wire                                        mgr35__std__lane15_strm1_data_valid  ,

            // manager 35, lane 16, stream 0      
            input   wire                                        std__mgr35__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane16_strm0_data        ,
            output  wire                                        mgr35__std__lane16_strm0_data_valid  ,

            // manager 35, lane 16, stream 1      
            input   wire                                        std__mgr35__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane16_strm1_data        ,
            output  wire                                        mgr35__std__lane16_strm1_data_valid  ,

            // manager 35, lane 17, stream 0      
            input   wire                                        std__mgr35__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane17_strm0_data        ,
            output  wire                                        mgr35__std__lane17_strm0_data_valid  ,

            // manager 35, lane 17, stream 1      
            input   wire                                        std__mgr35__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane17_strm1_data        ,
            output  wire                                        mgr35__std__lane17_strm1_data_valid  ,

            // manager 35, lane 18, stream 0      
            input   wire                                        std__mgr35__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane18_strm0_data        ,
            output  wire                                        mgr35__std__lane18_strm0_data_valid  ,

            // manager 35, lane 18, stream 1      
            input   wire                                        std__mgr35__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane18_strm1_data        ,
            output  wire                                        mgr35__std__lane18_strm1_data_valid  ,

            // manager 35, lane 19, stream 0      
            input   wire                                        std__mgr35__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane19_strm0_data        ,
            output  wire                                        mgr35__std__lane19_strm0_data_valid  ,

            // manager 35, lane 19, stream 1      
            input   wire                                        std__mgr35__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane19_strm1_data        ,
            output  wire                                        mgr35__std__lane19_strm1_data_valid  ,

            // manager 35, lane 20, stream 0      
            input   wire                                        std__mgr35__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane20_strm0_data        ,
            output  wire                                        mgr35__std__lane20_strm0_data_valid  ,

            // manager 35, lane 20, stream 1      
            input   wire                                        std__mgr35__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane20_strm1_data        ,
            output  wire                                        mgr35__std__lane20_strm1_data_valid  ,

            // manager 35, lane 21, stream 0      
            input   wire                                        std__mgr35__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane21_strm0_data        ,
            output  wire                                        mgr35__std__lane21_strm0_data_valid  ,

            // manager 35, lane 21, stream 1      
            input   wire                                        std__mgr35__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane21_strm1_data        ,
            output  wire                                        mgr35__std__lane21_strm1_data_valid  ,

            // manager 35, lane 22, stream 0      
            input   wire                                        std__mgr35__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane22_strm0_data        ,
            output  wire                                        mgr35__std__lane22_strm0_data_valid  ,

            // manager 35, lane 22, stream 1      
            input   wire                                        std__mgr35__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane22_strm1_data        ,
            output  wire                                        mgr35__std__lane22_strm1_data_valid  ,

            // manager 35, lane 23, stream 0      
            input   wire                                        std__mgr35__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane23_strm0_data        ,
            output  wire                                        mgr35__std__lane23_strm0_data_valid  ,

            // manager 35, lane 23, stream 1      
            input   wire                                        std__mgr35__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane23_strm1_data        ,
            output  wire                                        mgr35__std__lane23_strm1_data_valid  ,

            // manager 35, lane 24, stream 0      
            input   wire                                        std__mgr35__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane24_strm0_data        ,
            output  wire                                        mgr35__std__lane24_strm0_data_valid  ,

            // manager 35, lane 24, stream 1      
            input   wire                                        std__mgr35__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane24_strm1_data        ,
            output  wire                                        mgr35__std__lane24_strm1_data_valid  ,

            // manager 35, lane 25, stream 0      
            input   wire                                        std__mgr35__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane25_strm0_data        ,
            output  wire                                        mgr35__std__lane25_strm0_data_valid  ,

            // manager 35, lane 25, stream 1      
            input   wire                                        std__mgr35__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane25_strm1_data        ,
            output  wire                                        mgr35__std__lane25_strm1_data_valid  ,

            // manager 35, lane 26, stream 0      
            input   wire                                        std__mgr35__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane26_strm0_data        ,
            output  wire                                        mgr35__std__lane26_strm0_data_valid  ,

            // manager 35, lane 26, stream 1      
            input   wire                                        std__mgr35__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane26_strm1_data        ,
            output  wire                                        mgr35__std__lane26_strm1_data_valid  ,

            // manager 35, lane 27, stream 0      
            input   wire                                        std__mgr35__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane27_strm0_data        ,
            output  wire                                        mgr35__std__lane27_strm0_data_valid  ,

            // manager 35, lane 27, stream 1      
            input   wire                                        std__mgr35__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane27_strm1_data        ,
            output  wire                                        mgr35__std__lane27_strm1_data_valid  ,

            // manager 35, lane 28, stream 0      
            input   wire                                        std__mgr35__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane28_strm0_data        ,
            output  wire                                        mgr35__std__lane28_strm0_data_valid  ,

            // manager 35, lane 28, stream 1      
            input   wire                                        std__mgr35__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane28_strm1_data        ,
            output  wire                                        mgr35__std__lane28_strm1_data_valid  ,

            // manager 35, lane 29, stream 0      
            input   wire                                        std__mgr35__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane29_strm0_data        ,
            output  wire                                        mgr35__std__lane29_strm0_data_valid  ,

            // manager 35, lane 29, stream 1      
            input   wire                                        std__mgr35__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane29_strm1_data        ,
            output  wire                                        mgr35__std__lane29_strm1_data_valid  ,

            // manager 35, lane 30, stream 0      
            input   wire                                        std__mgr35__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane30_strm0_data        ,
            output  wire                                        mgr35__std__lane30_strm0_data_valid  ,

            // manager 35, lane 30, stream 1      
            input   wire                                        std__mgr35__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane30_strm1_data        ,
            output  wire                                        mgr35__std__lane30_strm1_data_valid  ,

            // manager 35, lane 31, stream 0      
            input   wire                                        std__mgr35__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane31_strm0_data        ,
            output  wire                                        mgr35__std__lane31_strm0_data_valid  ,

            // manager 35, lane 31, stream 1      
            input   wire                                        std__mgr35__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr35__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr35__std__lane31_strm1_data        ,
            output  wire                                        mgr35__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 36, lane 0, stream 0      
            input   wire                                        std__mgr36__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane0_strm0_data        ,
            output  wire                                        mgr36__std__lane0_strm0_data_valid  ,

            // manager 36, lane 0, stream 1      
            input   wire                                        std__mgr36__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane0_strm1_data        ,
            output  wire                                        mgr36__std__lane0_strm1_data_valid  ,

            // manager 36, lane 1, stream 0      
            input   wire                                        std__mgr36__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane1_strm0_data        ,
            output  wire                                        mgr36__std__lane1_strm0_data_valid  ,

            // manager 36, lane 1, stream 1      
            input   wire                                        std__mgr36__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane1_strm1_data        ,
            output  wire                                        mgr36__std__lane1_strm1_data_valid  ,

            // manager 36, lane 2, stream 0      
            input   wire                                        std__mgr36__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane2_strm0_data        ,
            output  wire                                        mgr36__std__lane2_strm0_data_valid  ,

            // manager 36, lane 2, stream 1      
            input   wire                                        std__mgr36__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane2_strm1_data        ,
            output  wire                                        mgr36__std__lane2_strm1_data_valid  ,

            // manager 36, lane 3, stream 0      
            input   wire                                        std__mgr36__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane3_strm0_data        ,
            output  wire                                        mgr36__std__lane3_strm0_data_valid  ,

            // manager 36, lane 3, stream 1      
            input   wire                                        std__mgr36__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane3_strm1_data        ,
            output  wire                                        mgr36__std__lane3_strm1_data_valid  ,

            // manager 36, lane 4, stream 0      
            input   wire                                        std__mgr36__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane4_strm0_data        ,
            output  wire                                        mgr36__std__lane4_strm0_data_valid  ,

            // manager 36, lane 4, stream 1      
            input   wire                                        std__mgr36__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane4_strm1_data        ,
            output  wire                                        mgr36__std__lane4_strm1_data_valid  ,

            // manager 36, lane 5, stream 0      
            input   wire                                        std__mgr36__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane5_strm0_data        ,
            output  wire                                        mgr36__std__lane5_strm0_data_valid  ,

            // manager 36, lane 5, stream 1      
            input   wire                                        std__mgr36__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane5_strm1_data        ,
            output  wire                                        mgr36__std__lane5_strm1_data_valid  ,

            // manager 36, lane 6, stream 0      
            input   wire                                        std__mgr36__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane6_strm0_data        ,
            output  wire                                        mgr36__std__lane6_strm0_data_valid  ,

            // manager 36, lane 6, stream 1      
            input   wire                                        std__mgr36__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane6_strm1_data        ,
            output  wire                                        mgr36__std__lane6_strm1_data_valid  ,

            // manager 36, lane 7, stream 0      
            input   wire                                        std__mgr36__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane7_strm0_data        ,
            output  wire                                        mgr36__std__lane7_strm0_data_valid  ,

            // manager 36, lane 7, stream 1      
            input   wire                                        std__mgr36__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane7_strm1_data        ,
            output  wire                                        mgr36__std__lane7_strm1_data_valid  ,

            // manager 36, lane 8, stream 0      
            input   wire                                        std__mgr36__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane8_strm0_data        ,
            output  wire                                        mgr36__std__lane8_strm0_data_valid  ,

            // manager 36, lane 8, stream 1      
            input   wire                                        std__mgr36__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane8_strm1_data        ,
            output  wire                                        mgr36__std__lane8_strm1_data_valid  ,

            // manager 36, lane 9, stream 0      
            input   wire                                        std__mgr36__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane9_strm0_data        ,
            output  wire                                        mgr36__std__lane9_strm0_data_valid  ,

            // manager 36, lane 9, stream 1      
            input   wire                                        std__mgr36__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane9_strm1_data        ,
            output  wire                                        mgr36__std__lane9_strm1_data_valid  ,

            // manager 36, lane 10, stream 0      
            input   wire                                        std__mgr36__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane10_strm0_data        ,
            output  wire                                        mgr36__std__lane10_strm0_data_valid  ,

            // manager 36, lane 10, stream 1      
            input   wire                                        std__mgr36__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane10_strm1_data        ,
            output  wire                                        mgr36__std__lane10_strm1_data_valid  ,

            // manager 36, lane 11, stream 0      
            input   wire                                        std__mgr36__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane11_strm0_data        ,
            output  wire                                        mgr36__std__lane11_strm0_data_valid  ,

            // manager 36, lane 11, stream 1      
            input   wire                                        std__mgr36__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane11_strm1_data        ,
            output  wire                                        mgr36__std__lane11_strm1_data_valid  ,

            // manager 36, lane 12, stream 0      
            input   wire                                        std__mgr36__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane12_strm0_data        ,
            output  wire                                        mgr36__std__lane12_strm0_data_valid  ,

            // manager 36, lane 12, stream 1      
            input   wire                                        std__mgr36__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane12_strm1_data        ,
            output  wire                                        mgr36__std__lane12_strm1_data_valid  ,

            // manager 36, lane 13, stream 0      
            input   wire                                        std__mgr36__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane13_strm0_data        ,
            output  wire                                        mgr36__std__lane13_strm0_data_valid  ,

            // manager 36, lane 13, stream 1      
            input   wire                                        std__mgr36__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane13_strm1_data        ,
            output  wire                                        mgr36__std__lane13_strm1_data_valid  ,

            // manager 36, lane 14, stream 0      
            input   wire                                        std__mgr36__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane14_strm0_data        ,
            output  wire                                        mgr36__std__lane14_strm0_data_valid  ,

            // manager 36, lane 14, stream 1      
            input   wire                                        std__mgr36__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane14_strm1_data        ,
            output  wire                                        mgr36__std__lane14_strm1_data_valid  ,

            // manager 36, lane 15, stream 0      
            input   wire                                        std__mgr36__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane15_strm0_data        ,
            output  wire                                        mgr36__std__lane15_strm0_data_valid  ,

            // manager 36, lane 15, stream 1      
            input   wire                                        std__mgr36__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane15_strm1_data        ,
            output  wire                                        mgr36__std__lane15_strm1_data_valid  ,

            // manager 36, lane 16, stream 0      
            input   wire                                        std__mgr36__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane16_strm0_data        ,
            output  wire                                        mgr36__std__lane16_strm0_data_valid  ,

            // manager 36, lane 16, stream 1      
            input   wire                                        std__mgr36__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane16_strm1_data        ,
            output  wire                                        mgr36__std__lane16_strm1_data_valid  ,

            // manager 36, lane 17, stream 0      
            input   wire                                        std__mgr36__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane17_strm0_data        ,
            output  wire                                        mgr36__std__lane17_strm0_data_valid  ,

            // manager 36, lane 17, stream 1      
            input   wire                                        std__mgr36__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane17_strm1_data        ,
            output  wire                                        mgr36__std__lane17_strm1_data_valid  ,

            // manager 36, lane 18, stream 0      
            input   wire                                        std__mgr36__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane18_strm0_data        ,
            output  wire                                        mgr36__std__lane18_strm0_data_valid  ,

            // manager 36, lane 18, stream 1      
            input   wire                                        std__mgr36__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane18_strm1_data        ,
            output  wire                                        mgr36__std__lane18_strm1_data_valid  ,

            // manager 36, lane 19, stream 0      
            input   wire                                        std__mgr36__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane19_strm0_data        ,
            output  wire                                        mgr36__std__lane19_strm0_data_valid  ,

            // manager 36, lane 19, stream 1      
            input   wire                                        std__mgr36__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane19_strm1_data        ,
            output  wire                                        mgr36__std__lane19_strm1_data_valid  ,

            // manager 36, lane 20, stream 0      
            input   wire                                        std__mgr36__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane20_strm0_data        ,
            output  wire                                        mgr36__std__lane20_strm0_data_valid  ,

            // manager 36, lane 20, stream 1      
            input   wire                                        std__mgr36__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane20_strm1_data        ,
            output  wire                                        mgr36__std__lane20_strm1_data_valid  ,

            // manager 36, lane 21, stream 0      
            input   wire                                        std__mgr36__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane21_strm0_data        ,
            output  wire                                        mgr36__std__lane21_strm0_data_valid  ,

            // manager 36, lane 21, stream 1      
            input   wire                                        std__mgr36__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane21_strm1_data        ,
            output  wire                                        mgr36__std__lane21_strm1_data_valid  ,

            // manager 36, lane 22, stream 0      
            input   wire                                        std__mgr36__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane22_strm0_data        ,
            output  wire                                        mgr36__std__lane22_strm0_data_valid  ,

            // manager 36, lane 22, stream 1      
            input   wire                                        std__mgr36__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane22_strm1_data        ,
            output  wire                                        mgr36__std__lane22_strm1_data_valid  ,

            // manager 36, lane 23, stream 0      
            input   wire                                        std__mgr36__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane23_strm0_data        ,
            output  wire                                        mgr36__std__lane23_strm0_data_valid  ,

            // manager 36, lane 23, stream 1      
            input   wire                                        std__mgr36__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane23_strm1_data        ,
            output  wire                                        mgr36__std__lane23_strm1_data_valid  ,

            // manager 36, lane 24, stream 0      
            input   wire                                        std__mgr36__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane24_strm0_data        ,
            output  wire                                        mgr36__std__lane24_strm0_data_valid  ,

            // manager 36, lane 24, stream 1      
            input   wire                                        std__mgr36__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane24_strm1_data        ,
            output  wire                                        mgr36__std__lane24_strm1_data_valid  ,

            // manager 36, lane 25, stream 0      
            input   wire                                        std__mgr36__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane25_strm0_data        ,
            output  wire                                        mgr36__std__lane25_strm0_data_valid  ,

            // manager 36, lane 25, stream 1      
            input   wire                                        std__mgr36__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane25_strm1_data        ,
            output  wire                                        mgr36__std__lane25_strm1_data_valid  ,

            // manager 36, lane 26, stream 0      
            input   wire                                        std__mgr36__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane26_strm0_data        ,
            output  wire                                        mgr36__std__lane26_strm0_data_valid  ,

            // manager 36, lane 26, stream 1      
            input   wire                                        std__mgr36__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane26_strm1_data        ,
            output  wire                                        mgr36__std__lane26_strm1_data_valid  ,

            // manager 36, lane 27, stream 0      
            input   wire                                        std__mgr36__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane27_strm0_data        ,
            output  wire                                        mgr36__std__lane27_strm0_data_valid  ,

            // manager 36, lane 27, stream 1      
            input   wire                                        std__mgr36__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane27_strm1_data        ,
            output  wire                                        mgr36__std__lane27_strm1_data_valid  ,

            // manager 36, lane 28, stream 0      
            input   wire                                        std__mgr36__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane28_strm0_data        ,
            output  wire                                        mgr36__std__lane28_strm0_data_valid  ,

            // manager 36, lane 28, stream 1      
            input   wire                                        std__mgr36__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane28_strm1_data        ,
            output  wire                                        mgr36__std__lane28_strm1_data_valid  ,

            // manager 36, lane 29, stream 0      
            input   wire                                        std__mgr36__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane29_strm0_data        ,
            output  wire                                        mgr36__std__lane29_strm0_data_valid  ,

            // manager 36, lane 29, stream 1      
            input   wire                                        std__mgr36__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane29_strm1_data        ,
            output  wire                                        mgr36__std__lane29_strm1_data_valid  ,

            // manager 36, lane 30, stream 0      
            input   wire                                        std__mgr36__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane30_strm0_data        ,
            output  wire                                        mgr36__std__lane30_strm0_data_valid  ,

            // manager 36, lane 30, stream 1      
            input   wire                                        std__mgr36__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane30_strm1_data        ,
            output  wire                                        mgr36__std__lane30_strm1_data_valid  ,

            // manager 36, lane 31, stream 0      
            input   wire                                        std__mgr36__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane31_strm0_data        ,
            output  wire                                        mgr36__std__lane31_strm0_data_valid  ,

            // manager 36, lane 31, stream 1      
            input   wire                                        std__mgr36__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr36__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr36__std__lane31_strm1_data        ,
            output  wire                                        mgr36__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 37, lane 0, stream 0      
            input   wire                                        std__mgr37__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane0_strm0_data        ,
            output  wire                                        mgr37__std__lane0_strm0_data_valid  ,

            // manager 37, lane 0, stream 1      
            input   wire                                        std__mgr37__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane0_strm1_data        ,
            output  wire                                        mgr37__std__lane0_strm1_data_valid  ,

            // manager 37, lane 1, stream 0      
            input   wire                                        std__mgr37__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane1_strm0_data        ,
            output  wire                                        mgr37__std__lane1_strm0_data_valid  ,

            // manager 37, lane 1, stream 1      
            input   wire                                        std__mgr37__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane1_strm1_data        ,
            output  wire                                        mgr37__std__lane1_strm1_data_valid  ,

            // manager 37, lane 2, stream 0      
            input   wire                                        std__mgr37__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane2_strm0_data        ,
            output  wire                                        mgr37__std__lane2_strm0_data_valid  ,

            // manager 37, lane 2, stream 1      
            input   wire                                        std__mgr37__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane2_strm1_data        ,
            output  wire                                        mgr37__std__lane2_strm1_data_valid  ,

            // manager 37, lane 3, stream 0      
            input   wire                                        std__mgr37__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane3_strm0_data        ,
            output  wire                                        mgr37__std__lane3_strm0_data_valid  ,

            // manager 37, lane 3, stream 1      
            input   wire                                        std__mgr37__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane3_strm1_data        ,
            output  wire                                        mgr37__std__lane3_strm1_data_valid  ,

            // manager 37, lane 4, stream 0      
            input   wire                                        std__mgr37__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane4_strm0_data        ,
            output  wire                                        mgr37__std__lane4_strm0_data_valid  ,

            // manager 37, lane 4, stream 1      
            input   wire                                        std__mgr37__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane4_strm1_data        ,
            output  wire                                        mgr37__std__lane4_strm1_data_valid  ,

            // manager 37, lane 5, stream 0      
            input   wire                                        std__mgr37__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane5_strm0_data        ,
            output  wire                                        mgr37__std__lane5_strm0_data_valid  ,

            // manager 37, lane 5, stream 1      
            input   wire                                        std__mgr37__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane5_strm1_data        ,
            output  wire                                        mgr37__std__lane5_strm1_data_valid  ,

            // manager 37, lane 6, stream 0      
            input   wire                                        std__mgr37__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane6_strm0_data        ,
            output  wire                                        mgr37__std__lane6_strm0_data_valid  ,

            // manager 37, lane 6, stream 1      
            input   wire                                        std__mgr37__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane6_strm1_data        ,
            output  wire                                        mgr37__std__lane6_strm1_data_valid  ,

            // manager 37, lane 7, stream 0      
            input   wire                                        std__mgr37__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane7_strm0_data        ,
            output  wire                                        mgr37__std__lane7_strm0_data_valid  ,

            // manager 37, lane 7, stream 1      
            input   wire                                        std__mgr37__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane7_strm1_data        ,
            output  wire                                        mgr37__std__lane7_strm1_data_valid  ,

            // manager 37, lane 8, stream 0      
            input   wire                                        std__mgr37__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane8_strm0_data        ,
            output  wire                                        mgr37__std__lane8_strm0_data_valid  ,

            // manager 37, lane 8, stream 1      
            input   wire                                        std__mgr37__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane8_strm1_data        ,
            output  wire                                        mgr37__std__lane8_strm1_data_valid  ,

            // manager 37, lane 9, stream 0      
            input   wire                                        std__mgr37__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane9_strm0_data        ,
            output  wire                                        mgr37__std__lane9_strm0_data_valid  ,

            // manager 37, lane 9, stream 1      
            input   wire                                        std__mgr37__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane9_strm1_data        ,
            output  wire                                        mgr37__std__lane9_strm1_data_valid  ,

            // manager 37, lane 10, stream 0      
            input   wire                                        std__mgr37__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane10_strm0_data        ,
            output  wire                                        mgr37__std__lane10_strm0_data_valid  ,

            // manager 37, lane 10, stream 1      
            input   wire                                        std__mgr37__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane10_strm1_data        ,
            output  wire                                        mgr37__std__lane10_strm1_data_valid  ,

            // manager 37, lane 11, stream 0      
            input   wire                                        std__mgr37__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane11_strm0_data        ,
            output  wire                                        mgr37__std__lane11_strm0_data_valid  ,

            // manager 37, lane 11, stream 1      
            input   wire                                        std__mgr37__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane11_strm1_data        ,
            output  wire                                        mgr37__std__lane11_strm1_data_valid  ,

            // manager 37, lane 12, stream 0      
            input   wire                                        std__mgr37__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane12_strm0_data        ,
            output  wire                                        mgr37__std__lane12_strm0_data_valid  ,

            // manager 37, lane 12, stream 1      
            input   wire                                        std__mgr37__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane12_strm1_data        ,
            output  wire                                        mgr37__std__lane12_strm1_data_valid  ,

            // manager 37, lane 13, stream 0      
            input   wire                                        std__mgr37__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane13_strm0_data        ,
            output  wire                                        mgr37__std__lane13_strm0_data_valid  ,

            // manager 37, lane 13, stream 1      
            input   wire                                        std__mgr37__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane13_strm1_data        ,
            output  wire                                        mgr37__std__lane13_strm1_data_valid  ,

            // manager 37, lane 14, stream 0      
            input   wire                                        std__mgr37__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane14_strm0_data        ,
            output  wire                                        mgr37__std__lane14_strm0_data_valid  ,

            // manager 37, lane 14, stream 1      
            input   wire                                        std__mgr37__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane14_strm1_data        ,
            output  wire                                        mgr37__std__lane14_strm1_data_valid  ,

            // manager 37, lane 15, stream 0      
            input   wire                                        std__mgr37__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane15_strm0_data        ,
            output  wire                                        mgr37__std__lane15_strm0_data_valid  ,

            // manager 37, lane 15, stream 1      
            input   wire                                        std__mgr37__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane15_strm1_data        ,
            output  wire                                        mgr37__std__lane15_strm1_data_valid  ,

            // manager 37, lane 16, stream 0      
            input   wire                                        std__mgr37__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane16_strm0_data        ,
            output  wire                                        mgr37__std__lane16_strm0_data_valid  ,

            // manager 37, lane 16, stream 1      
            input   wire                                        std__mgr37__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane16_strm1_data        ,
            output  wire                                        mgr37__std__lane16_strm1_data_valid  ,

            // manager 37, lane 17, stream 0      
            input   wire                                        std__mgr37__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane17_strm0_data        ,
            output  wire                                        mgr37__std__lane17_strm0_data_valid  ,

            // manager 37, lane 17, stream 1      
            input   wire                                        std__mgr37__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane17_strm1_data        ,
            output  wire                                        mgr37__std__lane17_strm1_data_valid  ,

            // manager 37, lane 18, stream 0      
            input   wire                                        std__mgr37__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane18_strm0_data        ,
            output  wire                                        mgr37__std__lane18_strm0_data_valid  ,

            // manager 37, lane 18, stream 1      
            input   wire                                        std__mgr37__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane18_strm1_data        ,
            output  wire                                        mgr37__std__lane18_strm1_data_valid  ,

            // manager 37, lane 19, stream 0      
            input   wire                                        std__mgr37__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane19_strm0_data        ,
            output  wire                                        mgr37__std__lane19_strm0_data_valid  ,

            // manager 37, lane 19, stream 1      
            input   wire                                        std__mgr37__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane19_strm1_data        ,
            output  wire                                        mgr37__std__lane19_strm1_data_valid  ,

            // manager 37, lane 20, stream 0      
            input   wire                                        std__mgr37__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane20_strm0_data        ,
            output  wire                                        mgr37__std__lane20_strm0_data_valid  ,

            // manager 37, lane 20, stream 1      
            input   wire                                        std__mgr37__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane20_strm1_data        ,
            output  wire                                        mgr37__std__lane20_strm1_data_valid  ,

            // manager 37, lane 21, stream 0      
            input   wire                                        std__mgr37__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane21_strm0_data        ,
            output  wire                                        mgr37__std__lane21_strm0_data_valid  ,

            // manager 37, lane 21, stream 1      
            input   wire                                        std__mgr37__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane21_strm1_data        ,
            output  wire                                        mgr37__std__lane21_strm1_data_valid  ,

            // manager 37, lane 22, stream 0      
            input   wire                                        std__mgr37__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane22_strm0_data        ,
            output  wire                                        mgr37__std__lane22_strm0_data_valid  ,

            // manager 37, lane 22, stream 1      
            input   wire                                        std__mgr37__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane22_strm1_data        ,
            output  wire                                        mgr37__std__lane22_strm1_data_valid  ,

            // manager 37, lane 23, stream 0      
            input   wire                                        std__mgr37__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane23_strm0_data        ,
            output  wire                                        mgr37__std__lane23_strm0_data_valid  ,

            // manager 37, lane 23, stream 1      
            input   wire                                        std__mgr37__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane23_strm1_data        ,
            output  wire                                        mgr37__std__lane23_strm1_data_valid  ,

            // manager 37, lane 24, stream 0      
            input   wire                                        std__mgr37__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane24_strm0_data        ,
            output  wire                                        mgr37__std__lane24_strm0_data_valid  ,

            // manager 37, lane 24, stream 1      
            input   wire                                        std__mgr37__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane24_strm1_data        ,
            output  wire                                        mgr37__std__lane24_strm1_data_valid  ,

            // manager 37, lane 25, stream 0      
            input   wire                                        std__mgr37__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane25_strm0_data        ,
            output  wire                                        mgr37__std__lane25_strm0_data_valid  ,

            // manager 37, lane 25, stream 1      
            input   wire                                        std__mgr37__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane25_strm1_data        ,
            output  wire                                        mgr37__std__lane25_strm1_data_valid  ,

            // manager 37, lane 26, stream 0      
            input   wire                                        std__mgr37__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane26_strm0_data        ,
            output  wire                                        mgr37__std__lane26_strm0_data_valid  ,

            // manager 37, lane 26, stream 1      
            input   wire                                        std__mgr37__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane26_strm1_data        ,
            output  wire                                        mgr37__std__lane26_strm1_data_valid  ,

            // manager 37, lane 27, stream 0      
            input   wire                                        std__mgr37__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane27_strm0_data        ,
            output  wire                                        mgr37__std__lane27_strm0_data_valid  ,

            // manager 37, lane 27, stream 1      
            input   wire                                        std__mgr37__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane27_strm1_data        ,
            output  wire                                        mgr37__std__lane27_strm1_data_valid  ,

            // manager 37, lane 28, stream 0      
            input   wire                                        std__mgr37__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane28_strm0_data        ,
            output  wire                                        mgr37__std__lane28_strm0_data_valid  ,

            // manager 37, lane 28, stream 1      
            input   wire                                        std__mgr37__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane28_strm1_data        ,
            output  wire                                        mgr37__std__lane28_strm1_data_valid  ,

            // manager 37, lane 29, stream 0      
            input   wire                                        std__mgr37__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane29_strm0_data        ,
            output  wire                                        mgr37__std__lane29_strm0_data_valid  ,

            // manager 37, lane 29, stream 1      
            input   wire                                        std__mgr37__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane29_strm1_data        ,
            output  wire                                        mgr37__std__lane29_strm1_data_valid  ,

            // manager 37, lane 30, stream 0      
            input   wire                                        std__mgr37__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane30_strm0_data        ,
            output  wire                                        mgr37__std__lane30_strm0_data_valid  ,

            // manager 37, lane 30, stream 1      
            input   wire                                        std__mgr37__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane30_strm1_data        ,
            output  wire                                        mgr37__std__lane30_strm1_data_valid  ,

            // manager 37, lane 31, stream 0      
            input   wire                                        std__mgr37__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane31_strm0_data        ,
            output  wire                                        mgr37__std__lane31_strm0_data_valid  ,

            // manager 37, lane 31, stream 1      
            input   wire                                        std__mgr37__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr37__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr37__std__lane31_strm1_data        ,
            output  wire                                        mgr37__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 38, lane 0, stream 0      
            input   wire                                        std__mgr38__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane0_strm0_data        ,
            output  wire                                        mgr38__std__lane0_strm0_data_valid  ,

            // manager 38, lane 0, stream 1      
            input   wire                                        std__mgr38__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane0_strm1_data        ,
            output  wire                                        mgr38__std__lane0_strm1_data_valid  ,

            // manager 38, lane 1, stream 0      
            input   wire                                        std__mgr38__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane1_strm0_data        ,
            output  wire                                        mgr38__std__lane1_strm0_data_valid  ,

            // manager 38, lane 1, stream 1      
            input   wire                                        std__mgr38__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane1_strm1_data        ,
            output  wire                                        mgr38__std__lane1_strm1_data_valid  ,

            // manager 38, lane 2, stream 0      
            input   wire                                        std__mgr38__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane2_strm0_data        ,
            output  wire                                        mgr38__std__lane2_strm0_data_valid  ,

            // manager 38, lane 2, stream 1      
            input   wire                                        std__mgr38__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane2_strm1_data        ,
            output  wire                                        mgr38__std__lane2_strm1_data_valid  ,

            // manager 38, lane 3, stream 0      
            input   wire                                        std__mgr38__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane3_strm0_data        ,
            output  wire                                        mgr38__std__lane3_strm0_data_valid  ,

            // manager 38, lane 3, stream 1      
            input   wire                                        std__mgr38__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane3_strm1_data        ,
            output  wire                                        mgr38__std__lane3_strm1_data_valid  ,

            // manager 38, lane 4, stream 0      
            input   wire                                        std__mgr38__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane4_strm0_data        ,
            output  wire                                        mgr38__std__lane4_strm0_data_valid  ,

            // manager 38, lane 4, stream 1      
            input   wire                                        std__mgr38__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane4_strm1_data        ,
            output  wire                                        mgr38__std__lane4_strm1_data_valid  ,

            // manager 38, lane 5, stream 0      
            input   wire                                        std__mgr38__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane5_strm0_data        ,
            output  wire                                        mgr38__std__lane5_strm0_data_valid  ,

            // manager 38, lane 5, stream 1      
            input   wire                                        std__mgr38__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane5_strm1_data        ,
            output  wire                                        mgr38__std__lane5_strm1_data_valid  ,

            // manager 38, lane 6, stream 0      
            input   wire                                        std__mgr38__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane6_strm0_data        ,
            output  wire                                        mgr38__std__lane6_strm0_data_valid  ,

            // manager 38, lane 6, stream 1      
            input   wire                                        std__mgr38__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane6_strm1_data        ,
            output  wire                                        mgr38__std__lane6_strm1_data_valid  ,

            // manager 38, lane 7, stream 0      
            input   wire                                        std__mgr38__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane7_strm0_data        ,
            output  wire                                        mgr38__std__lane7_strm0_data_valid  ,

            // manager 38, lane 7, stream 1      
            input   wire                                        std__mgr38__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane7_strm1_data        ,
            output  wire                                        mgr38__std__lane7_strm1_data_valid  ,

            // manager 38, lane 8, stream 0      
            input   wire                                        std__mgr38__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane8_strm0_data        ,
            output  wire                                        mgr38__std__lane8_strm0_data_valid  ,

            // manager 38, lane 8, stream 1      
            input   wire                                        std__mgr38__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane8_strm1_data        ,
            output  wire                                        mgr38__std__lane8_strm1_data_valid  ,

            // manager 38, lane 9, stream 0      
            input   wire                                        std__mgr38__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane9_strm0_data        ,
            output  wire                                        mgr38__std__lane9_strm0_data_valid  ,

            // manager 38, lane 9, stream 1      
            input   wire                                        std__mgr38__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane9_strm1_data        ,
            output  wire                                        mgr38__std__lane9_strm1_data_valid  ,

            // manager 38, lane 10, stream 0      
            input   wire                                        std__mgr38__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane10_strm0_data        ,
            output  wire                                        mgr38__std__lane10_strm0_data_valid  ,

            // manager 38, lane 10, stream 1      
            input   wire                                        std__mgr38__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane10_strm1_data        ,
            output  wire                                        mgr38__std__lane10_strm1_data_valid  ,

            // manager 38, lane 11, stream 0      
            input   wire                                        std__mgr38__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane11_strm0_data        ,
            output  wire                                        mgr38__std__lane11_strm0_data_valid  ,

            // manager 38, lane 11, stream 1      
            input   wire                                        std__mgr38__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane11_strm1_data        ,
            output  wire                                        mgr38__std__lane11_strm1_data_valid  ,

            // manager 38, lane 12, stream 0      
            input   wire                                        std__mgr38__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane12_strm0_data        ,
            output  wire                                        mgr38__std__lane12_strm0_data_valid  ,

            // manager 38, lane 12, stream 1      
            input   wire                                        std__mgr38__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane12_strm1_data        ,
            output  wire                                        mgr38__std__lane12_strm1_data_valid  ,

            // manager 38, lane 13, stream 0      
            input   wire                                        std__mgr38__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane13_strm0_data        ,
            output  wire                                        mgr38__std__lane13_strm0_data_valid  ,

            // manager 38, lane 13, stream 1      
            input   wire                                        std__mgr38__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane13_strm1_data        ,
            output  wire                                        mgr38__std__lane13_strm1_data_valid  ,

            // manager 38, lane 14, stream 0      
            input   wire                                        std__mgr38__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane14_strm0_data        ,
            output  wire                                        mgr38__std__lane14_strm0_data_valid  ,

            // manager 38, lane 14, stream 1      
            input   wire                                        std__mgr38__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane14_strm1_data        ,
            output  wire                                        mgr38__std__lane14_strm1_data_valid  ,

            // manager 38, lane 15, stream 0      
            input   wire                                        std__mgr38__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane15_strm0_data        ,
            output  wire                                        mgr38__std__lane15_strm0_data_valid  ,

            // manager 38, lane 15, stream 1      
            input   wire                                        std__mgr38__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane15_strm1_data        ,
            output  wire                                        mgr38__std__lane15_strm1_data_valid  ,

            // manager 38, lane 16, stream 0      
            input   wire                                        std__mgr38__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane16_strm0_data        ,
            output  wire                                        mgr38__std__lane16_strm0_data_valid  ,

            // manager 38, lane 16, stream 1      
            input   wire                                        std__mgr38__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane16_strm1_data        ,
            output  wire                                        mgr38__std__lane16_strm1_data_valid  ,

            // manager 38, lane 17, stream 0      
            input   wire                                        std__mgr38__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane17_strm0_data        ,
            output  wire                                        mgr38__std__lane17_strm0_data_valid  ,

            // manager 38, lane 17, stream 1      
            input   wire                                        std__mgr38__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane17_strm1_data        ,
            output  wire                                        mgr38__std__lane17_strm1_data_valid  ,

            // manager 38, lane 18, stream 0      
            input   wire                                        std__mgr38__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane18_strm0_data        ,
            output  wire                                        mgr38__std__lane18_strm0_data_valid  ,

            // manager 38, lane 18, stream 1      
            input   wire                                        std__mgr38__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane18_strm1_data        ,
            output  wire                                        mgr38__std__lane18_strm1_data_valid  ,

            // manager 38, lane 19, stream 0      
            input   wire                                        std__mgr38__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane19_strm0_data        ,
            output  wire                                        mgr38__std__lane19_strm0_data_valid  ,

            // manager 38, lane 19, stream 1      
            input   wire                                        std__mgr38__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane19_strm1_data        ,
            output  wire                                        mgr38__std__lane19_strm1_data_valid  ,

            // manager 38, lane 20, stream 0      
            input   wire                                        std__mgr38__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane20_strm0_data        ,
            output  wire                                        mgr38__std__lane20_strm0_data_valid  ,

            // manager 38, lane 20, stream 1      
            input   wire                                        std__mgr38__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane20_strm1_data        ,
            output  wire                                        mgr38__std__lane20_strm1_data_valid  ,

            // manager 38, lane 21, stream 0      
            input   wire                                        std__mgr38__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane21_strm0_data        ,
            output  wire                                        mgr38__std__lane21_strm0_data_valid  ,

            // manager 38, lane 21, stream 1      
            input   wire                                        std__mgr38__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane21_strm1_data        ,
            output  wire                                        mgr38__std__lane21_strm1_data_valid  ,

            // manager 38, lane 22, stream 0      
            input   wire                                        std__mgr38__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane22_strm0_data        ,
            output  wire                                        mgr38__std__lane22_strm0_data_valid  ,

            // manager 38, lane 22, stream 1      
            input   wire                                        std__mgr38__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane22_strm1_data        ,
            output  wire                                        mgr38__std__lane22_strm1_data_valid  ,

            // manager 38, lane 23, stream 0      
            input   wire                                        std__mgr38__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane23_strm0_data        ,
            output  wire                                        mgr38__std__lane23_strm0_data_valid  ,

            // manager 38, lane 23, stream 1      
            input   wire                                        std__mgr38__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane23_strm1_data        ,
            output  wire                                        mgr38__std__lane23_strm1_data_valid  ,

            // manager 38, lane 24, stream 0      
            input   wire                                        std__mgr38__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane24_strm0_data        ,
            output  wire                                        mgr38__std__lane24_strm0_data_valid  ,

            // manager 38, lane 24, stream 1      
            input   wire                                        std__mgr38__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane24_strm1_data        ,
            output  wire                                        mgr38__std__lane24_strm1_data_valid  ,

            // manager 38, lane 25, stream 0      
            input   wire                                        std__mgr38__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane25_strm0_data        ,
            output  wire                                        mgr38__std__lane25_strm0_data_valid  ,

            // manager 38, lane 25, stream 1      
            input   wire                                        std__mgr38__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane25_strm1_data        ,
            output  wire                                        mgr38__std__lane25_strm1_data_valid  ,

            // manager 38, lane 26, stream 0      
            input   wire                                        std__mgr38__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane26_strm0_data        ,
            output  wire                                        mgr38__std__lane26_strm0_data_valid  ,

            // manager 38, lane 26, stream 1      
            input   wire                                        std__mgr38__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane26_strm1_data        ,
            output  wire                                        mgr38__std__lane26_strm1_data_valid  ,

            // manager 38, lane 27, stream 0      
            input   wire                                        std__mgr38__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane27_strm0_data        ,
            output  wire                                        mgr38__std__lane27_strm0_data_valid  ,

            // manager 38, lane 27, stream 1      
            input   wire                                        std__mgr38__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane27_strm1_data        ,
            output  wire                                        mgr38__std__lane27_strm1_data_valid  ,

            // manager 38, lane 28, stream 0      
            input   wire                                        std__mgr38__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane28_strm0_data        ,
            output  wire                                        mgr38__std__lane28_strm0_data_valid  ,

            // manager 38, lane 28, stream 1      
            input   wire                                        std__mgr38__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane28_strm1_data        ,
            output  wire                                        mgr38__std__lane28_strm1_data_valid  ,

            // manager 38, lane 29, stream 0      
            input   wire                                        std__mgr38__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane29_strm0_data        ,
            output  wire                                        mgr38__std__lane29_strm0_data_valid  ,

            // manager 38, lane 29, stream 1      
            input   wire                                        std__mgr38__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane29_strm1_data        ,
            output  wire                                        mgr38__std__lane29_strm1_data_valid  ,

            // manager 38, lane 30, stream 0      
            input   wire                                        std__mgr38__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane30_strm0_data        ,
            output  wire                                        mgr38__std__lane30_strm0_data_valid  ,

            // manager 38, lane 30, stream 1      
            input   wire                                        std__mgr38__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane30_strm1_data        ,
            output  wire                                        mgr38__std__lane30_strm1_data_valid  ,

            // manager 38, lane 31, stream 0      
            input   wire                                        std__mgr38__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane31_strm0_data        ,
            output  wire                                        mgr38__std__lane31_strm0_data_valid  ,

            // manager 38, lane 31, stream 1      
            input   wire                                        std__mgr38__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr38__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr38__std__lane31_strm1_data        ,
            output  wire                                        mgr38__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 39, lane 0, stream 0      
            input   wire                                        std__mgr39__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane0_strm0_data        ,
            output  wire                                        mgr39__std__lane0_strm0_data_valid  ,

            // manager 39, lane 0, stream 1      
            input   wire                                        std__mgr39__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane0_strm1_data        ,
            output  wire                                        mgr39__std__lane0_strm1_data_valid  ,

            // manager 39, lane 1, stream 0      
            input   wire                                        std__mgr39__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane1_strm0_data        ,
            output  wire                                        mgr39__std__lane1_strm0_data_valid  ,

            // manager 39, lane 1, stream 1      
            input   wire                                        std__mgr39__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane1_strm1_data        ,
            output  wire                                        mgr39__std__lane1_strm1_data_valid  ,

            // manager 39, lane 2, stream 0      
            input   wire                                        std__mgr39__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane2_strm0_data        ,
            output  wire                                        mgr39__std__lane2_strm0_data_valid  ,

            // manager 39, lane 2, stream 1      
            input   wire                                        std__mgr39__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane2_strm1_data        ,
            output  wire                                        mgr39__std__lane2_strm1_data_valid  ,

            // manager 39, lane 3, stream 0      
            input   wire                                        std__mgr39__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane3_strm0_data        ,
            output  wire                                        mgr39__std__lane3_strm0_data_valid  ,

            // manager 39, lane 3, stream 1      
            input   wire                                        std__mgr39__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane3_strm1_data        ,
            output  wire                                        mgr39__std__lane3_strm1_data_valid  ,

            // manager 39, lane 4, stream 0      
            input   wire                                        std__mgr39__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane4_strm0_data        ,
            output  wire                                        mgr39__std__lane4_strm0_data_valid  ,

            // manager 39, lane 4, stream 1      
            input   wire                                        std__mgr39__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane4_strm1_data        ,
            output  wire                                        mgr39__std__lane4_strm1_data_valid  ,

            // manager 39, lane 5, stream 0      
            input   wire                                        std__mgr39__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane5_strm0_data        ,
            output  wire                                        mgr39__std__lane5_strm0_data_valid  ,

            // manager 39, lane 5, stream 1      
            input   wire                                        std__mgr39__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane5_strm1_data        ,
            output  wire                                        mgr39__std__lane5_strm1_data_valid  ,

            // manager 39, lane 6, stream 0      
            input   wire                                        std__mgr39__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane6_strm0_data        ,
            output  wire                                        mgr39__std__lane6_strm0_data_valid  ,

            // manager 39, lane 6, stream 1      
            input   wire                                        std__mgr39__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane6_strm1_data        ,
            output  wire                                        mgr39__std__lane6_strm1_data_valid  ,

            // manager 39, lane 7, stream 0      
            input   wire                                        std__mgr39__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane7_strm0_data        ,
            output  wire                                        mgr39__std__lane7_strm0_data_valid  ,

            // manager 39, lane 7, stream 1      
            input   wire                                        std__mgr39__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane7_strm1_data        ,
            output  wire                                        mgr39__std__lane7_strm1_data_valid  ,

            // manager 39, lane 8, stream 0      
            input   wire                                        std__mgr39__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane8_strm0_data        ,
            output  wire                                        mgr39__std__lane8_strm0_data_valid  ,

            // manager 39, lane 8, stream 1      
            input   wire                                        std__mgr39__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane8_strm1_data        ,
            output  wire                                        mgr39__std__lane8_strm1_data_valid  ,

            // manager 39, lane 9, stream 0      
            input   wire                                        std__mgr39__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane9_strm0_data        ,
            output  wire                                        mgr39__std__lane9_strm0_data_valid  ,

            // manager 39, lane 9, stream 1      
            input   wire                                        std__mgr39__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane9_strm1_data        ,
            output  wire                                        mgr39__std__lane9_strm1_data_valid  ,

            // manager 39, lane 10, stream 0      
            input   wire                                        std__mgr39__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane10_strm0_data        ,
            output  wire                                        mgr39__std__lane10_strm0_data_valid  ,

            // manager 39, lane 10, stream 1      
            input   wire                                        std__mgr39__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane10_strm1_data        ,
            output  wire                                        mgr39__std__lane10_strm1_data_valid  ,

            // manager 39, lane 11, stream 0      
            input   wire                                        std__mgr39__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane11_strm0_data        ,
            output  wire                                        mgr39__std__lane11_strm0_data_valid  ,

            // manager 39, lane 11, stream 1      
            input   wire                                        std__mgr39__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane11_strm1_data        ,
            output  wire                                        mgr39__std__lane11_strm1_data_valid  ,

            // manager 39, lane 12, stream 0      
            input   wire                                        std__mgr39__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane12_strm0_data        ,
            output  wire                                        mgr39__std__lane12_strm0_data_valid  ,

            // manager 39, lane 12, stream 1      
            input   wire                                        std__mgr39__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane12_strm1_data        ,
            output  wire                                        mgr39__std__lane12_strm1_data_valid  ,

            // manager 39, lane 13, stream 0      
            input   wire                                        std__mgr39__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane13_strm0_data        ,
            output  wire                                        mgr39__std__lane13_strm0_data_valid  ,

            // manager 39, lane 13, stream 1      
            input   wire                                        std__mgr39__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane13_strm1_data        ,
            output  wire                                        mgr39__std__lane13_strm1_data_valid  ,

            // manager 39, lane 14, stream 0      
            input   wire                                        std__mgr39__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane14_strm0_data        ,
            output  wire                                        mgr39__std__lane14_strm0_data_valid  ,

            // manager 39, lane 14, stream 1      
            input   wire                                        std__mgr39__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane14_strm1_data        ,
            output  wire                                        mgr39__std__lane14_strm1_data_valid  ,

            // manager 39, lane 15, stream 0      
            input   wire                                        std__mgr39__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane15_strm0_data        ,
            output  wire                                        mgr39__std__lane15_strm0_data_valid  ,

            // manager 39, lane 15, stream 1      
            input   wire                                        std__mgr39__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane15_strm1_data        ,
            output  wire                                        mgr39__std__lane15_strm1_data_valid  ,

            // manager 39, lane 16, stream 0      
            input   wire                                        std__mgr39__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane16_strm0_data        ,
            output  wire                                        mgr39__std__lane16_strm0_data_valid  ,

            // manager 39, lane 16, stream 1      
            input   wire                                        std__mgr39__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane16_strm1_data        ,
            output  wire                                        mgr39__std__lane16_strm1_data_valid  ,

            // manager 39, lane 17, stream 0      
            input   wire                                        std__mgr39__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane17_strm0_data        ,
            output  wire                                        mgr39__std__lane17_strm0_data_valid  ,

            // manager 39, lane 17, stream 1      
            input   wire                                        std__mgr39__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane17_strm1_data        ,
            output  wire                                        mgr39__std__lane17_strm1_data_valid  ,

            // manager 39, lane 18, stream 0      
            input   wire                                        std__mgr39__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane18_strm0_data        ,
            output  wire                                        mgr39__std__lane18_strm0_data_valid  ,

            // manager 39, lane 18, stream 1      
            input   wire                                        std__mgr39__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane18_strm1_data        ,
            output  wire                                        mgr39__std__lane18_strm1_data_valid  ,

            // manager 39, lane 19, stream 0      
            input   wire                                        std__mgr39__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane19_strm0_data        ,
            output  wire                                        mgr39__std__lane19_strm0_data_valid  ,

            // manager 39, lane 19, stream 1      
            input   wire                                        std__mgr39__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane19_strm1_data        ,
            output  wire                                        mgr39__std__lane19_strm1_data_valid  ,

            // manager 39, lane 20, stream 0      
            input   wire                                        std__mgr39__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane20_strm0_data        ,
            output  wire                                        mgr39__std__lane20_strm0_data_valid  ,

            // manager 39, lane 20, stream 1      
            input   wire                                        std__mgr39__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane20_strm1_data        ,
            output  wire                                        mgr39__std__lane20_strm1_data_valid  ,

            // manager 39, lane 21, stream 0      
            input   wire                                        std__mgr39__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane21_strm0_data        ,
            output  wire                                        mgr39__std__lane21_strm0_data_valid  ,

            // manager 39, lane 21, stream 1      
            input   wire                                        std__mgr39__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane21_strm1_data        ,
            output  wire                                        mgr39__std__lane21_strm1_data_valid  ,

            // manager 39, lane 22, stream 0      
            input   wire                                        std__mgr39__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane22_strm0_data        ,
            output  wire                                        mgr39__std__lane22_strm0_data_valid  ,

            // manager 39, lane 22, stream 1      
            input   wire                                        std__mgr39__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane22_strm1_data        ,
            output  wire                                        mgr39__std__lane22_strm1_data_valid  ,

            // manager 39, lane 23, stream 0      
            input   wire                                        std__mgr39__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane23_strm0_data        ,
            output  wire                                        mgr39__std__lane23_strm0_data_valid  ,

            // manager 39, lane 23, stream 1      
            input   wire                                        std__mgr39__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane23_strm1_data        ,
            output  wire                                        mgr39__std__lane23_strm1_data_valid  ,

            // manager 39, lane 24, stream 0      
            input   wire                                        std__mgr39__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane24_strm0_data        ,
            output  wire                                        mgr39__std__lane24_strm0_data_valid  ,

            // manager 39, lane 24, stream 1      
            input   wire                                        std__mgr39__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane24_strm1_data        ,
            output  wire                                        mgr39__std__lane24_strm1_data_valid  ,

            // manager 39, lane 25, stream 0      
            input   wire                                        std__mgr39__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane25_strm0_data        ,
            output  wire                                        mgr39__std__lane25_strm0_data_valid  ,

            // manager 39, lane 25, stream 1      
            input   wire                                        std__mgr39__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane25_strm1_data        ,
            output  wire                                        mgr39__std__lane25_strm1_data_valid  ,

            // manager 39, lane 26, stream 0      
            input   wire                                        std__mgr39__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane26_strm0_data        ,
            output  wire                                        mgr39__std__lane26_strm0_data_valid  ,

            // manager 39, lane 26, stream 1      
            input   wire                                        std__mgr39__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane26_strm1_data        ,
            output  wire                                        mgr39__std__lane26_strm1_data_valid  ,

            // manager 39, lane 27, stream 0      
            input   wire                                        std__mgr39__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane27_strm0_data        ,
            output  wire                                        mgr39__std__lane27_strm0_data_valid  ,

            // manager 39, lane 27, stream 1      
            input   wire                                        std__mgr39__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane27_strm1_data        ,
            output  wire                                        mgr39__std__lane27_strm1_data_valid  ,

            // manager 39, lane 28, stream 0      
            input   wire                                        std__mgr39__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane28_strm0_data        ,
            output  wire                                        mgr39__std__lane28_strm0_data_valid  ,

            // manager 39, lane 28, stream 1      
            input   wire                                        std__mgr39__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane28_strm1_data        ,
            output  wire                                        mgr39__std__lane28_strm1_data_valid  ,

            // manager 39, lane 29, stream 0      
            input   wire                                        std__mgr39__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane29_strm0_data        ,
            output  wire                                        mgr39__std__lane29_strm0_data_valid  ,

            // manager 39, lane 29, stream 1      
            input   wire                                        std__mgr39__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane29_strm1_data        ,
            output  wire                                        mgr39__std__lane29_strm1_data_valid  ,

            // manager 39, lane 30, stream 0      
            input   wire                                        std__mgr39__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane30_strm0_data        ,
            output  wire                                        mgr39__std__lane30_strm0_data_valid  ,

            // manager 39, lane 30, stream 1      
            input   wire                                        std__mgr39__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane30_strm1_data        ,
            output  wire                                        mgr39__std__lane30_strm1_data_valid  ,

            // manager 39, lane 31, stream 0      
            input   wire                                        std__mgr39__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane31_strm0_data        ,
            output  wire                                        mgr39__std__lane31_strm0_data_valid  ,

            // manager 39, lane 31, stream 1      
            input   wire                                        std__mgr39__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr39__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr39__std__lane31_strm1_data        ,
            output  wire                                        mgr39__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 40, lane 0, stream 0      
            input   wire                                        std__mgr40__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane0_strm0_data        ,
            output  wire                                        mgr40__std__lane0_strm0_data_valid  ,

            // manager 40, lane 0, stream 1      
            input   wire                                        std__mgr40__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane0_strm1_data        ,
            output  wire                                        mgr40__std__lane0_strm1_data_valid  ,

            // manager 40, lane 1, stream 0      
            input   wire                                        std__mgr40__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane1_strm0_data        ,
            output  wire                                        mgr40__std__lane1_strm0_data_valid  ,

            // manager 40, lane 1, stream 1      
            input   wire                                        std__mgr40__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane1_strm1_data        ,
            output  wire                                        mgr40__std__lane1_strm1_data_valid  ,

            // manager 40, lane 2, stream 0      
            input   wire                                        std__mgr40__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane2_strm0_data        ,
            output  wire                                        mgr40__std__lane2_strm0_data_valid  ,

            // manager 40, lane 2, stream 1      
            input   wire                                        std__mgr40__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane2_strm1_data        ,
            output  wire                                        mgr40__std__lane2_strm1_data_valid  ,

            // manager 40, lane 3, stream 0      
            input   wire                                        std__mgr40__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane3_strm0_data        ,
            output  wire                                        mgr40__std__lane3_strm0_data_valid  ,

            // manager 40, lane 3, stream 1      
            input   wire                                        std__mgr40__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane3_strm1_data        ,
            output  wire                                        mgr40__std__lane3_strm1_data_valid  ,

            // manager 40, lane 4, stream 0      
            input   wire                                        std__mgr40__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane4_strm0_data        ,
            output  wire                                        mgr40__std__lane4_strm0_data_valid  ,

            // manager 40, lane 4, stream 1      
            input   wire                                        std__mgr40__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane4_strm1_data        ,
            output  wire                                        mgr40__std__lane4_strm1_data_valid  ,

            // manager 40, lane 5, stream 0      
            input   wire                                        std__mgr40__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane5_strm0_data        ,
            output  wire                                        mgr40__std__lane5_strm0_data_valid  ,

            // manager 40, lane 5, stream 1      
            input   wire                                        std__mgr40__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane5_strm1_data        ,
            output  wire                                        mgr40__std__lane5_strm1_data_valid  ,

            // manager 40, lane 6, stream 0      
            input   wire                                        std__mgr40__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane6_strm0_data        ,
            output  wire                                        mgr40__std__lane6_strm0_data_valid  ,

            // manager 40, lane 6, stream 1      
            input   wire                                        std__mgr40__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane6_strm1_data        ,
            output  wire                                        mgr40__std__lane6_strm1_data_valid  ,

            // manager 40, lane 7, stream 0      
            input   wire                                        std__mgr40__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane7_strm0_data        ,
            output  wire                                        mgr40__std__lane7_strm0_data_valid  ,

            // manager 40, lane 7, stream 1      
            input   wire                                        std__mgr40__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane7_strm1_data        ,
            output  wire                                        mgr40__std__lane7_strm1_data_valid  ,

            // manager 40, lane 8, stream 0      
            input   wire                                        std__mgr40__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane8_strm0_data        ,
            output  wire                                        mgr40__std__lane8_strm0_data_valid  ,

            // manager 40, lane 8, stream 1      
            input   wire                                        std__mgr40__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane8_strm1_data        ,
            output  wire                                        mgr40__std__lane8_strm1_data_valid  ,

            // manager 40, lane 9, stream 0      
            input   wire                                        std__mgr40__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane9_strm0_data        ,
            output  wire                                        mgr40__std__lane9_strm0_data_valid  ,

            // manager 40, lane 9, stream 1      
            input   wire                                        std__mgr40__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane9_strm1_data        ,
            output  wire                                        mgr40__std__lane9_strm1_data_valid  ,

            // manager 40, lane 10, stream 0      
            input   wire                                        std__mgr40__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane10_strm0_data        ,
            output  wire                                        mgr40__std__lane10_strm0_data_valid  ,

            // manager 40, lane 10, stream 1      
            input   wire                                        std__mgr40__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane10_strm1_data        ,
            output  wire                                        mgr40__std__lane10_strm1_data_valid  ,

            // manager 40, lane 11, stream 0      
            input   wire                                        std__mgr40__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane11_strm0_data        ,
            output  wire                                        mgr40__std__lane11_strm0_data_valid  ,

            // manager 40, lane 11, stream 1      
            input   wire                                        std__mgr40__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane11_strm1_data        ,
            output  wire                                        mgr40__std__lane11_strm1_data_valid  ,

            // manager 40, lane 12, stream 0      
            input   wire                                        std__mgr40__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane12_strm0_data        ,
            output  wire                                        mgr40__std__lane12_strm0_data_valid  ,

            // manager 40, lane 12, stream 1      
            input   wire                                        std__mgr40__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane12_strm1_data        ,
            output  wire                                        mgr40__std__lane12_strm1_data_valid  ,

            // manager 40, lane 13, stream 0      
            input   wire                                        std__mgr40__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane13_strm0_data        ,
            output  wire                                        mgr40__std__lane13_strm0_data_valid  ,

            // manager 40, lane 13, stream 1      
            input   wire                                        std__mgr40__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane13_strm1_data        ,
            output  wire                                        mgr40__std__lane13_strm1_data_valid  ,

            // manager 40, lane 14, stream 0      
            input   wire                                        std__mgr40__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane14_strm0_data        ,
            output  wire                                        mgr40__std__lane14_strm0_data_valid  ,

            // manager 40, lane 14, stream 1      
            input   wire                                        std__mgr40__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane14_strm1_data        ,
            output  wire                                        mgr40__std__lane14_strm1_data_valid  ,

            // manager 40, lane 15, stream 0      
            input   wire                                        std__mgr40__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane15_strm0_data        ,
            output  wire                                        mgr40__std__lane15_strm0_data_valid  ,

            // manager 40, lane 15, stream 1      
            input   wire                                        std__mgr40__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane15_strm1_data        ,
            output  wire                                        mgr40__std__lane15_strm1_data_valid  ,

            // manager 40, lane 16, stream 0      
            input   wire                                        std__mgr40__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane16_strm0_data        ,
            output  wire                                        mgr40__std__lane16_strm0_data_valid  ,

            // manager 40, lane 16, stream 1      
            input   wire                                        std__mgr40__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane16_strm1_data        ,
            output  wire                                        mgr40__std__lane16_strm1_data_valid  ,

            // manager 40, lane 17, stream 0      
            input   wire                                        std__mgr40__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane17_strm0_data        ,
            output  wire                                        mgr40__std__lane17_strm0_data_valid  ,

            // manager 40, lane 17, stream 1      
            input   wire                                        std__mgr40__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane17_strm1_data        ,
            output  wire                                        mgr40__std__lane17_strm1_data_valid  ,

            // manager 40, lane 18, stream 0      
            input   wire                                        std__mgr40__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane18_strm0_data        ,
            output  wire                                        mgr40__std__lane18_strm0_data_valid  ,

            // manager 40, lane 18, stream 1      
            input   wire                                        std__mgr40__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane18_strm1_data        ,
            output  wire                                        mgr40__std__lane18_strm1_data_valid  ,

            // manager 40, lane 19, stream 0      
            input   wire                                        std__mgr40__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane19_strm0_data        ,
            output  wire                                        mgr40__std__lane19_strm0_data_valid  ,

            // manager 40, lane 19, stream 1      
            input   wire                                        std__mgr40__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane19_strm1_data        ,
            output  wire                                        mgr40__std__lane19_strm1_data_valid  ,

            // manager 40, lane 20, stream 0      
            input   wire                                        std__mgr40__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane20_strm0_data        ,
            output  wire                                        mgr40__std__lane20_strm0_data_valid  ,

            // manager 40, lane 20, stream 1      
            input   wire                                        std__mgr40__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane20_strm1_data        ,
            output  wire                                        mgr40__std__lane20_strm1_data_valid  ,

            // manager 40, lane 21, stream 0      
            input   wire                                        std__mgr40__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane21_strm0_data        ,
            output  wire                                        mgr40__std__lane21_strm0_data_valid  ,

            // manager 40, lane 21, stream 1      
            input   wire                                        std__mgr40__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane21_strm1_data        ,
            output  wire                                        mgr40__std__lane21_strm1_data_valid  ,

            // manager 40, lane 22, stream 0      
            input   wire                                        std__mgr40__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane22_strm0_data        ,
            output  wire                                        mgr40__std__lane22_strm0_data_valid  ,

            // manager 40, lane 22, stream 1      
            input   wire                                        std__mgr40__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane22_strm1_data        ,
            output  wire                                        mgr40__std__lane22_strm1_data_valid  ,

            // manager 40, lane 23, stream 0      
            input   wire                                        std__mgr40__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane23_strm0_data        ,
            output  wire                                        mgr40__std__lane23_strm0_data_valid  ,

            // manager 40, lane 23, stream 1      
            input   wire                                        std__mgr40__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane23_strm1_data        ,
            output  wire                                        mgr40__std__lane23_strm1_data_valid  ,

            // manager 40, lane 24, stream 0      
            input   wire                                        std__mgr40__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane24_strm0_data        ,
            output  wire                                        mgr40__std__lane24_strm0_data_valid  ,

            // manager 40, lane 24, stream 1      
            input   wire                                        std__mgr40__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane24_strm1_data        ,
            output  wire                                        mgr40__std__lane24_strm1_data_valid  ,

            // manager 40, lane 25, stream 0      
            input   wire                                        std__mgr40__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane25_strm0_data        ,
            output  wire                                        mgr40__std__lane25_strm0_data_valid  ,

            // manager 40, lane 25, stream 1      
            input   wire                                        std__mgr40__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane25_strm1_data        ,
            output  wire                                        mgr40__std__lane25_strm1_data_valid  ,

            // manager 40, lane 26, stream 0      
            input   wire                                        std__mgr40__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane26_strm0_data        ,
            output  wire                                        mgr40__std__lane26_strm0_data_valid  ,

            // manager 40, lane 26, stream 1      
            input   wire                                        std__mgr40__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane26_strm1_data        ,
            output  wire                                        mgr40__std__lane26_strm1_data_valid  ,

            // manager 40, lane 27, stream 0      
            input   wire                                        std__mgr40__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane27_strm0_data        ,
            output  wire                                        mgr40__std__lane27_strm0_data_valid  ,

            // manager 40, lane 27, stream 1      
            input   wire                                        std__mgr40__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane27_strm1_data        ,
            output  wire                                        mgr40__std__lane27_strm1_data_valid  ,

            // manager 40, lane 28, stream 0      
            input   wire                                        std__mgr40__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane28_strm0_data        ,
            output  wire                                        mgr40__std__lane28_strm0_data_valid  ,

            // manager 40, lane 28, stream 1      
            input   wire                                        std__mgr40__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane28_strm1_data        ,
            output  wire                                        mgr40__std__lane28_strm1_data_valid  ,

            // manager 40, lane 29, stream 0      
            input   wire                                        std__mgr40__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane29_strm0_data        ,
            output  wire                                        mgr40__std__lane29_strm0_data_valid  ,

            // manager 40, lane 29, stream 1      
            input   wire                                        std__mgr40__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane29_strm1_data        ,
            output  wire                                        mgr40__std__lane29_strm1_data_valid  ,

            // manager 40, lane 30, stream 0      
            input   wire                                        std__mgr40__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane30_strm0_data        ,
            output  wire                                        mgr40__std__lane30_strm0_data_valid  ,

            // manager 40, lane 30, stream 1      
            input   wire                                        std__mgr40__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane30_strm1_data        ,
            output  wire                                        mgr40__std__lane30_strm1_data_valid  ,

            // manager 40, lane 31, stream 0      
            input   wire                                        std__mgr40__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane31_strm0_data        ,
            output  wire                                        mgr40__std__lane31_strm0_data_valid  ,

            // manager 40, lane 31, stream 1      
            input   wire                                        std__mgr40__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr40__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr40__std__lane31_strm1_data        ,
            output  wire                                        mgr40__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 41, lane 0, stream 0      
            input   wire                                        std__mgr41__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane0_strm0_data        ,
            output  wire                                        mgr41__std__lane0_strm0_data_valid  ,

            // manager 41, lane 0, stream 1      
            input   wire                                        std__mgr41__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane0_strm1_data        ,
            output  wire                                        mgr41__std__lane0_strm1_data_valid  ,

            // manager 41, lane 1, stream 0      
            input   wire                                        std__mgr41__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane1_strm0_data        ,
            output  wire                                        mgr41__std__lane1_strm0_data_valid  ,

            // manager 41, lane 1, stream 1      
            input   wire                                        std__mgr41__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane1_strm1_data        ,
            output  wire                                        mgr41__std__lane1_strm1_data_valid  ,

            // manager 41, lane 2, stream 0      
            input   wire                                        std__mgr41__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane2_strm0_data        ,
            output  wire                                        mgr41__std__lane2_strm0_data_valid  ,

            // manager 41, lane 2, stream 1      
            input   wire                                        std__mgr41__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane2_strm1_data        ,
            output  wire                                        mgr41__std__lane2_strm1_data_valid  ,

            // manager 41, lane 3, stream 0      
            input   wire                                        std__mgr41__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane3_strm0_data        ,
            output  wire                                        mgr41__std__lane3_strm0_data_valid  ,

            // manager 41, lane 3, stream 1      
            input   wire                                        std__mgr41__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane3_strm1_data        ,
            output  wire                                        mgr41__std__lane3_strm1_data_valid  ,

            // manager 41, lane 4, stream 0      
            input   wire                                        std__mgr41__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane4_strm0_data        ,
            output  wire                                        mgr41__std__lane4_strm0_data_valid  ,

            // manager 41, lane 4, stream 1      
            input   wire                                        std__mgr41__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane4_strm1_data        ,
            output  wire                                        mgr41__std__lane4_strm1_data_valid  ,

            // manager 41, lane 5, stream 0      
            input   wire                                        std__mgr41__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane5_strm0_data        ,
            output  wire                                        mgr41__std__lane5_strm0_data_valid  ,

            // manager 41, lane 5, stream 1      
            input   wire                                        std__mgr41__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane5_strm1_data        ,
            output  wire                                        mgr41__std__lane5_strm1_data_valid  ,

            // manager 41, lane 6, stream 0      
            input   wire                                        std__mgr41__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane6_strm0_data        ,
            output  wire                                        mgr41__std__lane6_strm0_data_valid  ,

            // manager 41, lane 6, stream 1      
            input   wire                                        std__mgr41__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane6_strm1_data        ,
            output  wire                                        mgr41__std__lane6_strm1_data_valid  ,

            // manager 41, lane 7, stream 0      
            input   wire                                        std__mgr41__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane7_strm0_data        ,
            output  wire                                        mgr41__std__lane7_strm0_data_valid  ,

            // manager 41, lane 7, stream 1      
            input   wire                                        std__mgr41__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane7_strm1_data        ,
            output  wire                                        mgr41__std__lane7_strm1_data_valid  ,

            // manager 41, lane 8, stream 0      
            input   wire                                        std__mgr41__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane8_strm0_data        ,
            output  wire                                        mgr41__std__lane8_strm0_data_valid  ,

            // manager 41, lane 8, stream 1      
            input   wire                                        std__mgr41__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane8_strm1_data        ,
            output  wire                                        mgr41__std__lane8_strm1_data_valid  ,

            // manager 41, lane 9, stream 0      
            input   wire                                        std__mgr41__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane9_strm0_data        ,
            output  wire                                        mgr41__std__lane9_strm0_data_valid  ,

            // manager 41, lane 9, stream 1      
            input   wire                                        std__mgr41__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane9_strm1_data        ,
            output  wire                                        mgr41__std__lane9_strm1_data_valid  ,

            // manager 41, lane 10, stream 0      
            input   wire                                        std__mgr41__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane10_strm0_data        ,
            output  wire                                        mgr41__std__lane10_strm0_data_valid  ,

            // manager 41, lane 10, stream 1      
            input   wire                                        std__mgr41__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane10_strm1_data        ,
            output  wire                                        mgr41__std__lane10_strm1_data_valid  ,

            // manager 41, lane 11, stream 0      
            input   wire                                        std__mgr41__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane11_strm0_data        ,
            output  wire                                        mgr41__std__lane11_strm0_data_valid  ,

            // manager 41, lane 11, stream 1      
            input   wire                                        std__mgr41__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane11_strm1_data        ,
            output  wire                                        mgr41__std__lane11_strm1_data_valid  ,

            // manager 41, lane 12, stream 0      
            input   wire                                        std__mgr41__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane12_strm0_data        ,
            output  wire                                        mgr41__std__lane12_strm0_data_valid  ,

            // manager 41, lane 12, stream 1      
            input   wire                                        std__mgr41__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane12_strm1_data        ,
            output  wire                                        mgr41__std__lane12_strm1_data_valid  ,

            // manager 41, lane 13, stream 0      
            input   wire                                        std__mgr41__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane13_strm0_data        ,
            output  wire                                        mgr41__std__lane13_strm0_data_valid  ,

            // manager 41, lane 13, stream 1      
            input   wire                                        std__mgr41__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane13_strm1_data        ,
            output  wire                                        mgr41__std__lane13_strm1_data_valid  ,

            // manager 41, lane 14, stream 0      
            input   wire                                        std__mgr41__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane14_strm0_data        ,
            output  wire                                        mgr41__std__lane14_strm0_data_valid  ,

            // manager 41, lane 14, stream 1      
            input   wire                                        std__mgr41__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane14_strm1_data        ,
            output  wire                                        mgr41__std__lane14_strm1_data_valid  ,

            // manager 41, lane 15, stream 0      
            input   wire                                        std__mgr41__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane15_strm0_data        ,
            output  wire                                        mgr41__std__lane15_strm0_data_valid  ,

            // manager 41, lane 15, stream 1      
            input   wire                                        std__mgr41__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane15_strm1_data        ,
            output  wire                                        mgr41__std__lane15_strm1_data_valid  ,

            // manager 41, lane 16, stream 0      
            input   wire                                        std__mgr41__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane16_strm0_data        ,
            output  wire                                        mgr41__std__lane16_strm0_data_valid  ,

            // manager 41, lane 16, stream 1      
            input   wire                                        std__mgr41__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane16_strm1_data        ,
            output  wire                                        mgr41__std__lane16_strm1_data_valid  ,

            // manager 41, lane 17, stream 0      
            input   wire                                        std__mgr41__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane17_strm0_data        ,
            output  wire                                        mgr41__std__lane17_strm0_data_valid  ,

            // manager 41, lane 17, stream 1      
            input   wire                                        std__mgr41__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane17_strm1_data        ,
            output  wire                                        mgr41__std__lane17_strm1_data_valid  ,

            // manager 41, lane 18, stream 0      
            input   wire                                        std__mgr41__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane18_strm0_data        ,
            output  wire                                        mgr41__std__lane18_strm0_data_valid  ,

            // manager 41, lane 18, stream 1      
            input   wire                                        std__mgr41__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane18_strm1_data        ,
            output  wire                                        mgr41__std__lane18_strm1_data_valid  ,

            // manager 41, lane 19, stream 0      
            input   wire                                        std__mgr41__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane19_strm0_data        ,
            output  wire                                        mgr41__std__lane19_strm0_data_valid  ,

            // manager 41, lane 19, stream 1      
            input   wire                                        std__mgr41__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane19_strm1_data        ,
            output  wire                                        mgr41__std__lane19_strm1_data_valid  ,

            // manager 41, lane 20, stream 0      
            input   wire                                        std__mgr41__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane20_strm0_data        ,
            output  wire                                        mgr41__std__lane20_strm0_data_valid  ,

            // manager 41, lane 20, stream 1      
            input   wire                                        std__mgr41__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane20_strm1_data        ,
            output  wire                                        mgr41__std__lane20_strm1_data_valid  ,

            // manager 41, lane 21, stream 0      
            input   wire                                        std__mgr41__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane21_strm0_data        ,
            output  wire                                        mgr41__std__lane21_strm0_data_valid  ,

            // manager 41, lane 21, stream 1      
            input   wire                                        std__mgr41__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane21_strm1_data        ,
            output  wire                                        mgr41__std__lane21_strm1_data_valid  ,

            // manager 41, lane 22, stream 0      
            input   wire                                        std__mgr41__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane22_strm0_data        ,
            output  wire                                        mgr41__std__lane22_strm0_data_valid  ,

            // manager 41, lane 22, stream 1      
            input   wire                                        std__mgr41__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane22_strm1_data        ,
            output  wire                                        mgr41__std__lane22_strm1_data_valid  ,

            // manager 41, lane 23, stream 0      
            input   wire                                        std__mgr41__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane23_strm0_data        ,
            output  wire                                        mgr41__std__lane23_strm0_data_valid  ,

            // manager 41, lane 23, stream 1      
            input   wire                                        std__mgr41__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane23_strm1_data        ,
            output  wire                                        mgr41__std__lane23_strm1_data_valid  ,

            // manager 41, lane 24, stream 0      
            input   wire                                        std__mgr41__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane24_strm0_data        ,
            output  wire                                        mgr41__std__lane24_strm0_data_valid  ,

            // manager 41, lane 24, stream 1      
            input   wire                                        std__mgr41__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane24_strm1_data        ,
            output  wire                                        mgr41__std__lane24_strm1_data_valid  ,

            // manager 41, lane 25, stream 0      
            input   wire                                        std__mgr41__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane25_strm0_data        ,
            output  wire                                        mgr41__std__lane25_strm0_data_valid  ,

            // manager 41, lane 25, stream 1      
            input   wire                                        std__mgr41__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane25_strm1_data        ,
            output  wire                                        mgr41__std__lane25_strm1_data_valid  ,

            // manager 41, lane 26, stream 0      
            input   wire                                        std__mgr41__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane26_strm0_data        ,
            output  wire                                        mgr41__std__lane26_strm0_data_valid  ,

            // manager 41, lane 26, stream 1      
            input   wire                                        std__mgr41__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane26_strm1_data        ,
            output  wire                                        mgr41__std__lane26_strm1_data_valid  ,

            // manager 41, lane 27, stream 0      
            input   wire                                        std__mgr41__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane27_strm0_data        ,
            output  wire                                        mgr41__std__lane27_strm0_data_valid  ,

            // manager 41, lane 27, stream 1      
            input   wire                                        std__mgr41__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane27_strm1_data        ,
            output  wire                                        mgr41__std__lane27_strm1_data_valid  ,

            // manager 41, lane 28, stream 0      
            input   wire                                        std__mgr41__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane28_strm0_data        ,
            output  wire                                        mgr41__std__lane28_strm0_data_valid  ,

            // manager 41, lane 28, stream 1      
            input   wire                                        std__mgr41__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane28_strm1_data        ,
            output  wire                                        mgr41__std__lane28_strm1_data_valid  ,

            // manager 41, lane 29, stream 0      
            input   wire                                        std__mgr41__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane29_strm0_data        ,
            output  wire                                        mgr41__std__lane29_strm0_data_valid  ,

            // manager 41, lane 29, stream 1      
            input   wire                                        std__mgr41__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane29_strm1_data        ,
            output  wire                                        mgr41__std__lane29_strm1_data_valid  ,

            // manager 41, lane 30, stream 0      
            input   wire                                        std__mgr41__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane30_strm0_data        ,
            output  wire                                        mgr41__std__lane30_strm0_data_valid  ,

            // manager 41, lane 30, stream 1      
            input   wire                                        std__mgr41__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane30_strm1_data        ,
            output  wire                                        mgr41__std__lane30_strm1_data_valid  ,

            // manager 41, lane 31, stream 0      
            input   wire                                        std__mgr41__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane31_strm0_data        ,
            output  wire                                        mgr41__std__lane31_strm0_data_valid  ,

            // manager 41, lane 31, stream 1      
            input   wire                                        std__mgr41__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr41__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr41__std__lane31_strm1_data        ,
            output  wire                                        mgr41__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 42, lane 0, stream 0      
            input   wire                                        std__mgr42__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane0_strm0_data        ,
            output  wire                                        mgr42__std__lane0_strm0_data_valid  ,

            // manager 42, lane 0, stream 1      
            input   wire                                        std__mgr42__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane0_strm1_data        ,
            output  wire                                        mgr42__std__lane0_strm1_data_valid  ,

            // manager 42, lane 1, stream 0      
            input   wire                                        std__mgr42__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane1_strm0_data        ,
            output  wire                                        mgr42__std__lane1_strm0_data_valid  ,

            // manager 42, lane 1, stream 1      
            input   wire                                        std__mgr42__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane1_strm1_data        ,
            output  wire                                        mgr42__std__lane1_strm1_data_valid  ,

            // manager 42, lane 2, stream 0      
            input   wire                                        std__mgr42__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane2_strm0_data        ,
            output  wire                                        mgr42__std__lane2_strm0_data_valid  ,

            // manager 42, lane 2, stream 1      
            input   wire                                        std__mgr42__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane2_strm1_data        ,
            output  wire                                        mgr42__std__lane2_strm1_data_valid  ,

            // manager 42, lane 3, stream 0      
            input   wire                                        std__mgr42__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane3_strm0_data        ,
            output  wire                                        mgr42__std__lane3_strm0_data_valid  ,

            // manager 42, lane 3, stream 1      
            input   wire                                        std__mgr42__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane3_strm1_data        ,
            output  wire                                        mgr42__std__lane3_strm1_data_valid  ,

            // manager 42, lane 4, stream 0      
            input   wire                                        std__mgr42__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane4_strm0_data        ,
            output  wire                                        mgr42__std__lane4_strm0_data_valid  ,

            // manager 42, lane 4, stream 1      
            input   wire                                        std__mgr42__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane4_strm1_data        ,
            output  wire                                        mgr42__std__lane4_strm1_data_valid  ,

            // manager 42, lane 5, stream 0      
            input   wire                                        std__mgr42__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane5_strm0_data        ,
            output  wire                                        mgr42__std__lane5_strm0_data_valid  ,

            // manager 42, lane 5, stream 1      
            input   wire                                        std__mgr42__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane5_strm1_data        ,
            output  wire                                        mgr42__std__lane5_strm1_data_valid  ,

            // manager 42, lane 6, stream 0      
            input   wire                                        std__mgr42__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane6_strm0_data        ,
            output  wire                                        mgr42__std__lane6_strm0_data_valid  ,

            // manager 42, lane 6, stream 1      
            input   wire                                        std__mgr42__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane6_strm1_data        ,
            output  wire                                        mgr42__std__lane6_strm1_data_valid  ,

            // manager 42, lane 7, stream 0      
            input   wire                                        std__mgr42__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane7_strm0_data        ,
            output  wire                                        mgr42__std__lane7_strm0_data_valid  ,

            // manager 42, lane 7, stream 1      
            input   wire                                        std__mgr42__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane7_strm1_data        ,
            output  wire                                        mgr42__std__lane7_strm1_data_valid  ,

            // manager 42, lane 8, stream 0      
            input   wire                                        std__mgr42__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane8_strm0_data        ,
            output  wire                                        mgr42__std__lane8_strm0_data_valid  ,

            // manager 42, lane 8, stream 1      
            input   wire                                        std__mgr42__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane8_strm1_data        ,
            output  wire                                        mgr42__std__lane8_strm1_data_valid  ,

            // manager 42, lane 9, stream 0      
            input   wire                                        std__mgr42__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane9_strm0_data        ,
            output  wire                                        mgr42__std__lane9_strm0_data_valid  ,

            // manager 42, lane 9, stream 1      
            input   wire                                        std__mgr42__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane9_strm1_data        ,
            output  wire                                        mgr42__std__lane9_strm1_data_valid  ,

            // manager 42, lane 10, stream 0      
            input   wire                                        std__mgr42__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane10_strm0_data        ,
            output  wire                                        mgr42__std__lane10_strm0_data_valid  ,

            // manager 42, lane 10, stream 1      
            input   wire                                        std__mgr42__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane10_strm1_data        ,
            output  wire                                        mgr42__std__lane10_strm1_data_valid  ,

            // manager 42, lane 11, stream 0      
            input   wire                                        std__mgr42__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane11_strm0_data        ,
            output  wire                                        mgr42__std__lane11_strm0_data_valid  ,

            // manager 42, lane 11, stream 1      
            input   wire                                        std__mgr42__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane11_strm1_data        ,
            output  wire                                        mgr42__std__lane11_strm1_data_valid  ,

            // manager 42, lane 12, stream 0      
            input   wire                                        std__mgr42__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane12_strm0_data        ,
            output  wire                                        mgr42__std__lane12_strm0_data_valid  ,

            // manager 42, lane 12, stream 1      
            input   wire                                        std__mgr42__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane12_strm1_data        ,
            output  wire                                        mgr42__std__lane12_strm1_data_valid  ,

            // manager 42, lane 13, stream 0      
            input   wire                                        std__mgr42__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane13_strm0_data        ,
            output  wire                                        mgr42__std__lane13_strm0_data_valid  ,

            // manager 42, lane 13, stream 1      
            input   wire                                        std__mgr42__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane13_strm1_data        ,
            output  wire                                        mgr42__std__lane13_strm1_data_valid  ,

            // manager 42, lane 14, stream 0      
            input   wire                                        std__mgr42__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane14_strm0_data        ,
            output  wire                                        mgr42__std__lane14_strm0_data_valid  ,

            // manager 42, lane 14, stream 1      
            input   wire                                        std__mgr42__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane14_strm1_data        ,
            output  wire                                        mgr42__std__lane14_strm1_data_valid  ,

            // manager 42, lane 15, stream 0      
            input   wire                                        std__mgr42__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane15_strm0_data        ,
            output  wire                                        mgr42__std__lane15_strm0_data_valid  ,

            // manager 42, lane 15, stream 1      
            input   wire                                        std__mgr42__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane15_strm1_data        ,
            output  wire                                        mgr42__std__lane15_strm1_data_valid  ,

            // manager 42, lane 16, stream 0      
            input   wire                                        std__mgr42__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane16_strm0_data        ,
            output  wire                                        mgr42__std__lane16_strm0_data_valid  ,

            // manager 42, lane 16, stream 1      
            input   wire                                        std__mgr42__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane16_strm1_data        ,
            output  wire                                        mgr42__std__lane16_strm1_data_valid  ,

            // manager 42, lane 17, stream 0      
            input   wire                                        std__mgr42__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane17_strm0_data        ,
            output  wire                                        mgr42__std__lane17_strm0_data_valid  ,

            // manager 42, lane 17, stream 1      
            input   wire                                        std__mgr42__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane17_strm1_data        ,
            output  wire                                        mgr42__std__lane17_strm1_data_valid  ,

            // manager 42, lane 18, stream 0      
            input   wire                                        std__mgr42__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane18_strm0_data        ,
            output  wire                                        mgr42__std__lane18_strm0_data_valid  ,

            // manager 42, lane 18, stream 1      
            input   wire                                        std__mgr42__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane18_strm1_data        ,
            output  wire                                        mgr42__std__lane18_strm1_data_valid  ,

            // manager 42, lane 19, stream 0      
            input   wire                                        std__mgr42__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane19_strm0_data        ,
            output  wire                                        mgr42__std__lane19_strm0_data_valid  ,

            // manager 42, lane 19, stream 1      
            input   wire                                        std__mgr42__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane19_strm1_data        ,
            output  wire                                        mgr42__std__lane19_strm1_data_valid  ,

            // manager 42, lane 20, stream 0      
            input   wire                                        std__mgr42__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane20_strm0_data        ,
            output  wire                                        mgr42__std__lane20_strm0_data_valid  ,

            // manager 42, lane 20, stream 1      
            input   wire                                        std__mgr42__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane20_strm1_data        ,
            output  wire                                        mgr42__std__lane20_strm1_data_valid  ,

            // manager 42, lane 21, stream 0      
            input   wire                                        std__mgr42__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane21_strm0_data        ,
            output  wire                                        mgr42__std__lane21_strm0_data_valid  ,

            // manager 42, lane 21, stream 1      
            input   wire                                        std__mgr42__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane21_strm1_data        ,
            output  wire                                        mgr42__std__lane21_strm1_data_valid  ,

            // manager 42, lane 22, stream 0      
            input   wire                                        std__mgr42__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane22_strm0_data        ,
            output  wire                                        mgr42__std__lane22_strm0_data_valid  ,

            // manager 42, lane 22, stream 1      
            input   wire                                        std__mgr42__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane22_strm1_data        ,
            output  wire                                        mgr42__std__lane22_strm1_data_valid  ,

            // manager 42, lane 23, stream 0      
            input   wire                                        std__mgr42__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane23_strm0_data        ,
            output  wire                                        mgr42__std__lane23_strm0_data_valid  ,

            // manager 42, lane 23, stream 1      
            input   wire                                        std__mgr42__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane23_strm1_data        ,
            output  wire                                        mgr42__std__lane23_strm1_data_valid  ,

            // manager 42, lane 24, stream 0      
            input   wire                                        std__mgr42__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane24_strm0_data        ,
            output  wire                                        mgr42__std__lane24_strm0_data_valid  ,

            // manager 42, lane 24, stream 1      
            input   wire                                        std__mgr42__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane24_strm1_data        ,
            output  wire                                        mgr42__std__lane24_strm1_data_valid  ,

            // manager 42, lane 25, stream 0      
            input   wire                                        std__mgr42__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane25_strm0_data        ,
            output  wire                                        mgr42__std__lane25_strm0_data_valid  ,

            // manager 42, lane 25, stream 1      
            input   wire                                        std__mgr42__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane25_strm1_data        ,
            output  wire                                        mgr42__std__lane25_strm1_data_valid  ,

            // manager 42, lane 26, stream 0      
            input   wire                                        std__mgr42__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane26_strm0_data        ,
            output  wire                                        mgr42__std__lane26_strm0_data_valid  ,

            // manager 42, lane 26, stream 1      
            input   wire                                        std__mgr42__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane26_strm1_data        ,
            output  wire                                        mgr42__std__lane26_strm1_data_valid  ,

            // manager 42, lane 27, stream 0      
            input   wire                                        std__mgr42__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane27_strm0_data        ,
            output  wire                                        mgr42__std__lane27_strm0_data_valid  ,

            // manager 42, lane 27, stream 1      
            input   wire                                        std__mgr42__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane27_strm1_data        ,
            output  wire                                        mgr42__std__lane27_strm1_data_valid  ,

            // manager 42, lane 28, stream 0      
            input   wire                                        std__mgr42__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane28_strm0_data        ,
            output  wire                                        mgr42__std__lane28_strm0_data_valid  ,

            // manager 42, lane 28, stream 1      
            input   wire                                        std__mgr42__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane28_strm1_data        ,
            output  wire                                        mgr42__std__lane28_strm1_data_valid  ,

            // manager 42, lane 29, stream 0      
            input   wire                                        std__mgr42__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane29_strm0_data        ,
            output  wire                                        mgr42__std__lane29_strm0_data_valid  ,

            // manager 42, lane 29, stream 1      
            input   wire                                        std__mgr42__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane29_strm1_data        ,
            output  wire                                        mgr42__std__lane29_strm1_data_valid  ,

            // manager 42, lane 30, stream 0      
            input   wire                                        std__mgr42__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane30_strm0_data        ,
            output  wire                                        mgr42__std__lane30_strm0_data_valid  ,

            // manager 42, lane 30, stream 1      
            input   wire                                        std__mgr42__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane30_strm1_data        ,
            output  wire                                        mgr42__std__lane30_strm1_data_valid  ,

            // manager 42, lane 31, stream 0      
            input   wire                                        std__mgr42__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane31_strm0_data        ,
            output  wire                                        mgr42__std__lane31_strm0_data_valid  ,

            // manager 42, lane 31, stream 1      
            input   wire                                        std__mgr42__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr42__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr42__std__lane31_strm1_data        ,
            output  wire                                        mgr42__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 43, lane 0, stream 0      
            input   wire                                        std__mgr43__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane0_strm0_data        ,
            output  wire                                        mgr43__std__lane0_strm0_data_valid  ,

            // manager 43, lane 0, stream 1      
            input   wire                                        std__mgr43__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane0_strm1_data        ,
            output  wire                                        mgr43__std__lane0_strm1_data_valid  ,

            // manager 43, lane 1, stream 0      
            input   wire                                        std__mgr43__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane1_strm0_data        ,
            output  wire                                        mgr43__std__lane1_strm0_data_valid  ,

            // manager 43, lane 1, stream 1      
            input   wire                                        std__mgr43__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane1_strm1_data        ,
            output  wire                                        mgr43__std__lane1_strm1_data_valid  ,

            // manager 43, lane 2, stream 0      
            input   wire                                        std__mgr43__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane2_strm0_data        ,
            output  wire                                        mgr43__std__lane2_strm0_data_valid  ,

            // manager 43, lane 2, stream 1      
            input   wire                                        std__mgr43__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane2_strm1_data        ,
            output  wire                                        mgr43__std__lane2_strm1_data_valid  ,

            // manager 43, lane 3, stream 0      
            input   wire                                        std__mgr43__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane3_strm0_data        ,
            output  wire                                        mgr43__std__lane3_strm0_data_valid  ,

            // manager 43, lane 3, stream 1      
            input   wire                                        std__mgr43__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane3_strm1_data        ,
            output  wire                                        mgr43__std__lane3_strm1_data_valid  ,

            // manager 43, lane 4, stream 0      
            input   wire                                        std__mgr43__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane4_strm0_data        ,
            output  wire                                        mgr43__std__lane4_strm0_data_valid  ,

            // manager 43, lane 4, stream 1      
            input   wire                                        std__mgr43__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane4_strm1_data        ,
            output  wire                                        mgr43__std__lane4_strm1_data_valid  ,

            // manager 43, lane 5, stream 0      
            input   wire                                        std__mgr43__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane5_strm0_data        ,
            output  wire                                        mgr43__std__lane5_strm0_data_valid  ,

            // manager 43, lane 5, stream 1      
            input   wire                                        std__mgr43__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane5_strm1_data        ,
            output  wire                                        mgr43__std__lane5_strm1_data_valid  ,

            // manager 43, lane 6, stream 0      
            input   wire                                        std__mgr43__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane6_strm0_data        ,
            output  wire                                        mgr43__std__lane6_strm0_data_valid  ,

            // manager 43, lane 6, stream 1      
            input   wire                                        std__mgr43__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane6_strm1_data        ,
            output  wire                                        mgr43__std__lane6_strm1_data_valid  ,

            // manager 43, lane 7, stream 0      
            input   wire                                        std__mgr43__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane7_strm0_data        ,
            output  wire                                        mgr43__std__lane7_strm0_data_valid  ,

            // manager 43, lane 7, stream 1      
            input   wire                                        std__mgr43__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane7_strm1_data        ,
            output  wire                                        mgr43__std__lane7_strm1_data_valid  ,

            // manager 43, lane 8, stream 0      
            input   wire                                        std__mgr43__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane8_strm0_data        ,
            output  wire                                        mgr43__std__lane8_strm0_data_valid  ,

            // manager 43, lane 8, stream 1      
            input   wire                                        std__mgr43__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane8_strm1_data        ,
            output  wire                                        mgr43__std__lane8_strm1_data_valid  ,

            // manager 43, lane 9, stream 0      
            input   wire                                        std__mgr43__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane9_strm0_data        ,
            output  wire                                        mgr43__std__lane9_strm0_data_valid  ,

            // manager 43, lane 9, stream 1      
            input   wire                                        std__mgr43__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane9_strm1_data        ,
            output  wire                                        mgr43__std__lane9_strm1_data_valid  ,

            // manager 43, lane 10, stream 0      
            input   wire                                        std__mgr43__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane10_strm0_data        ,
            output  wire                                        mgr43__std__lane10_strm0_data_valid  ,

            // manager 43, lane 10, stream 1      
            input   wire                                        std__mgr43__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane10_strm1_data        ,
            output  wire                                        mgr43__std__lane10_strm1_data_valid  ,

            // manager 43, lane 11, stream 0      
            input   wire                                        std__mgr43__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane11_strm0_data        ,
            output  wire                                        mgr43__std__lane11_strm0_data_valid  ,

            // manager 43, lane 11, stream 1      
            input   wire                                        std__mgr43__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane11_strm1_data        ,
            output  wire                                        mgr43__std__lane11_strm1_data_valid  ,

            // manager 43, lane 12, stream 0      
            input   wire                                        std__mgr43__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane12_strm0_data        ,
            output  wire                                        mgr43__std__lane12_strm0_data_valid  ,

            // manager 43, lane 12, stream 1      
            input   wire                                        std__mgr43__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane12_strm1_data        ,
            output  wire                                        mgr43__std__lane12_strm1_data_valid  ,

            // manager 43, lane 13, stream 0      
            input   wire                                        std__mgr43__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane13_strm0_data        ,
            output  wire                                        mgr43__std__lane13_strm0_data_valid  ,

            // manager 43, lane 13, stream 1      
            input   wire                                        std__mgr43__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane13_strm1_data        ,
            output  wire                                        mgr43__std__lane13_strm1_data_valid  ,

            // manager 43, lane 14, stream 0      
            input   wire                                        std__mgr43__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane14_strm0_data        ,
            output  wire                                        mgr43__std__lane14_strm0_data_valid  ,

            // manager 43, lane 14, stream 1      
            input   wire                                        std__mgr43__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane14_strm1_data        ,
            output  wire                                        mgr43__std__lane14_strm1_data_valid  ,

            // manager 43, lane 15, stream 0      
            input   wire                                        std__mgr43__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane15_strm0_data        ,
            output  wire                                        mgr43__std__lane15_strm0_data_valid  ,

            // manager 43, lane 15, stream 1      
            input   wire                                        std__mgr43__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane15_strm1_data        ,
            output  wire                                        mgr43__std__lane15_strm1_data_valid  ,

            // manager 43, lane 16, stream 0      
            input   wire                                        std__mgr43__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane16_strm0_data        ,
            output  wire                                        mgr43__std__lane16_strm0_data_valid  ,

            // manager 43, lane 16, stream 1      
            input   wire                                        std__mgr43__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane16_strm1_data        ,
            output  wire                                        mgr43__std__lane16_strm1_data_valid  ,

            // manager 43, lane 17, stream 0      
            input   wire                                        std__mgr43__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane17_strm0_data        ,
            output  wire                                        mgr43__std__lane17_strm0_data_valid  ,

            // manager 43, lane 17, stream 1      
            input   wire                                        std__mgr43__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane17_strm1_data        ,
            output  wire                                        mgr43__std__lane17_strm1_data_valid  ,

            // manager 43, lane 18, stream 0      
            input   wire                                        std__mgr43__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane18_strm0_data        ,
            output  wire                                        mgr43__std__lane18_strm0_data_valid  ,

            // manager 43, lane 18, stream 1      
            input   wire                                        std__mgr43__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane18_strm1_data        ,
            output  wire                                        mgr43__std__lane18_strm1_data_valid  ,

            // manager 43, lane 19, stream 0      
            input   wire                                        std__mgr43__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane19_strm0_data        ,
            output  wire                                        mgr43__std__lane19_strm0_data_valid  ,

            // manager 43, lane 19, stream 1      
            input   wire                                        std__mgr43__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane19_strm1_data        ,
            output  wire                                        mgr43__std__lane19_strm1_data_valid  ,

            // manager 43, lane 20, stream 0      
            input   wire                                        std__mgr43__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane20_strm0_data        ,
            output  wire                                        mgr43__std__lane20_strm0_data_valid  ,

            // manager 43, lane 20, stream 1      
            input   wire                                        std__mgr43__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane20_strm1_data        ,
            output  wire                                        mgr43__std__lane20_strm1_data_valid  ,

            // manager 43, lane 21, stream 0      
            input   wire                                        std__mgr43__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane21_strm0_data        ,
            output  wire                                        mgr43__std__lane21_strm0_data_valid  ,

            // manager 43, lane 21, stream 1      
            input   wire                                        std__mgr43__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane21_strm1_data        ,
            output  wire                                        mgr43__std__lane21_strm1_data_valid  ,

            // manager 43, lane 22, stream 0      
            input   wire                                        std__mgr43__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane22_strm0_data        ,
            output  wire                                        mgr43__std__lane22_strm0_data_valid  ,

            // manager 43, lane 22, stream 1      
            input   wire                                        std__mgr43__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane22_strm1_data        ,
            output  wire                                        mgr43__std__lane22_strm1_data_valid  ,

            // manager 43, lane 23, stream 0      
            input   wire                                        std__mgr43__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane23_strm0_data        ,
            output  wire                                        mgr43__std__lane23_strm0_data_valid  ,

            // manager 43, lane 23, stream 1      
            input   wire                                        std__mgr43__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane23_strm1_data        ,
            output  wire                                        mgr43__std__lane23_strm1_data_valid  ,

            // manager 43, lane 24, stream 0      
            input   wire                                        std__mgr43__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane24_strm0_data        ,
            output  wire                                        mgr43__std__lane24_strm0_data_valid  ,

            // manager 43, lane 24, stream 1      
            input   wire                                        std__mgr43__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane24_strm1_data        ,
            output  wire                                        mgr43__std__lane24_strm1_data_valid  ,

            // manager 43, lane 25, stream 0      
            input   wire                                        std__mgr43__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane25_strm0_data        ,
            output  wire                                        mgr43__std__lane25_strm0_data_valid  ,

            // manager 43, lane 25, stream 1      
            input   wire                                        std__mgr43__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane25_strm1_data        ,
            output  wire                                        mgr43__std__lane25_strm1_data_valid  ,

            // manager 43, lane 26, stream 0      
            input   wire                                        std__mgr43__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane26_strm0_data        ,
            output  wire                                        mgr43__std__lane26_strm0_data_valid  ,

            // manager 43, lane 26, stream 1      
            input   wire                                        std__mgr43__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane26_strm1_data        ,
            output  wire                                        mgr43__std__lane26_strm1_data_valid  ,

            // manager 43, lane 27, stream 0      
            input   wire                                        std__mgr43__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane27_strm0_data        ,
            output  wire                                        mgr43__std__lane27_strm0_data_valid  ,

            // manager 43, lane 27, stream 1      
            input   wire                                        std__mgr43__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane27_strm1_data        ,
            output  wire                                        mgr43__std__lane27_strm1_data_valid  ,

            // manager 43, lane 28, stream 0      
            input   wire                                        std__mgr43__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane28_strm0_data        ,
            output  wire                                        mgr43__std__lane28_strm0_data_valid  ,

            // manager 43, lane 28, stream 1      
            input   wire                                        std__mgr43__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane28_strm1_data        ,
            output  wire                                        mgr43__std__lane28_strm1_data_valid  ,

            // manager 43, lane 29, stream 0      
            input   wire                                        std__mgr43__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane29_strm0_data        ,
            output  wire                                        mgr43__std__lane29_strm0_data_valid  ,

            // manager 43, lane 29, stream 1      
            input   wire                                        std__mgr43__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane29_strm1_data        ,
            output  wire                                        mgr43__std__lane29_strm1_data_valid  ,

            // manager 43, lane 30, stream 0      
            input   wire                                        std__mgr43__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane30_strm0_data        ,
            output  wire                                        mgr43__std__lane30_strm0_data_valid  ,

            // manager 43, lane 30, stream 1      
            input   wire                                        std__mgr43__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane30_strm1_data        ,
            output  wire                                        mgr43__std__lane30_strm1_data_valid  ,

            // manager 43, lane 31, stream 0      
            input   wire                                        std__mgr43__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane31_strm0_data        ,
            output  wire                                        mgr43__std__lane31_strm0_data_valid  ,

            // manager 43, lane 31, stream 1      
            input   wire                                        std__mgr43__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr43__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr43__std__lane31_strm1_data        ,
            output  wire                                        mgr43__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 44, lane 0, stream 0      
            input   wire                                        std__mgr44__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane0_strm0_data        ,
            output  wire                                        mgr44__std__lane0_strm0_data_valid  ,

            // manager 44, lane 0, stream 1      
            input   wire                                        std__mgr44__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane0_strm1_data        ,
            output  wire                                        mgr44__std__lane0_strm1_data_valid  ,

            // manager 44, lane 1, stream 0      
            input   wire                                        std__mgr44__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane1_strm0_data        ,
            output  wire                                        mgr44__std__lane1_strm0_data_valid  ,

            // manager 44, lane 1, stream 1      
            input   wire                                        std__mgr44__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane1_strm1_data        ,
            output  wire                                        mgr44__std__lane1_strm1_data_valid  ,

            // manager 44, lane 2, stream 0      
            input   wire                                        std__mgr44__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane2_strm0_data        ,
            output  wire                                        mgr44__std__lane2_strm0_data_valid  ,

            // manager 44, lane 2, stream 1      
            input   wire                                        std__mgr44__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane2_strm1_data        ,
            output  wire                                        mgr44__std__lane2_strm1_data_valid  ,

            // manager 44, lane 3, stream 0      
            input   wire                                        std__mgr44__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane3_strm0_data        ,
            output  wire                                        mgr44__std__lane3_strm0_data_valid  ,

            // manager 44, lane 3, stream 1      
            input   wire                                        std__mgr44__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane3_strm1_data        ,
            output  wire                                        mgr44__std__lane3_strm1_data_valid  ,

            // manager 44, lane 4, stream 0      
            input   wire                                        std__mgr44__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane4_strm0_data        ,
            output  wire                                        mgr44__std__lane4_strm0_data_valid  ,

            // manager 44, lane 4, stream 1      
            input   wire                                        std__mgr44__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane4_strm1_data        ,
            output  wire                                        mgr44__std__lane4_strm1_data_valid  ,

            // manager 44, lane 5, stream 0      
            input   wire                                        std__mgr44__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane5_strm0_data        ,
            output  wire                                        mgr44__std__lane5_strm0_data_valid  ,

            // manager 44, lane 5, stream 1      
            input   wire                                        std__mgr44__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane5_strm1_data        ,
            output  wire                                        mgr44__std__lane5_strm1_data_valid  ,

            // manager 44, lane 6, stream 0      
            input   wire                                        std__mgr44__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane6_strm0_data        ,
            output  wire                                        mgr44__std__lane6_strm0_data_valid  ,

            // manager 44, lane 6, stream 1      
            input   wire                                        std__mgr44__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane6_strm1_data        ,
            output  wire                                        mgr44__std__lane6_strm1_data_valid  ,

            // manager 44, lane 7, stream 0      
            input   wire                                        std__mgr44__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane7_strm0_data        ,
            output  wire                                        mgr44__std__lane7_strm0_data_valid  ,

            // manager 44, lane 7, stream 1      
            input   wire                                        std__mgr44__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane7_strm1_data        ,
            output  wire                                        mgr44__std__lane7_strm1_data_valid  ,

            // manager 44, lane 8, stream 0      
            input   wire                                        std__mgr44__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane8_strm0_data        ,
            output  wire                                        mgr44__std__lane8_strm0_data_valid  ,

            // manager 44, lane 8, stream 1      
            input   wire                                        std__mgr44__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane8_strm1_data        ,
            output  wire                                        mgr44__std__lane8_strm1_data_valid  ,

            // manager 44, lane 9, stream 0      
            input   wire                                        std__mgr44__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane9_strm0_data        ,
            output  wire                                        mgr44__std__lane9_strm0_data_valid  ,

            // manager 44, lane 9, stream 1      
            input   wire                                        std__mgr44__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane9_strm1_data        ,
            output  wire                                        mgr44__std__lane9_strm1_data_valid  ,

            // manager 44, lane 10, stream 0      
            input   wire                                        std__mgr44__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane10_strm0_data        ,
            output  wire                                        mgr44__std__lane10_strm0_data_valid  ,

            // manager 44, lane 10, stream 1      
            input   wire                                        std__mgr44__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane10_strm1_data        ,
            output  wire                                        mgr44__std__lane10_strm1_data_valid  ,

            // manager 44, lane 11, stream 0      
            input   wire                                        std__mgr44__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane11_strm0_data        ,
            output  wire                                        mgr44__std__lane11_strm0_data_valid  ,

            // manager 44, lane 11, stream 1      
            input   wire                                        std__mgr44__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane11_strm1_data        ,
            output  wire                                        mgr44__std__lane11_strm1_data_valid  ,

            // manager 44, lane 12, stream 0      
            input   wire                                        std__mgr44__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane12_strm0_data        ,
            output  wire                                        mgr44__std__lane12_strm0_data_valid  ,

            // manager 44, lane 12, stream 1      
            input   wire                                        std__mgr44__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane12_strm1_data        ,
            output  wire                                        mgr44__std__lane12_strm1_data_valid  ,

            // manager 44, lane 13, stream 0      
            input   wire                                        std__mgr44__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane13_strm0_data        ,
            output  wire                                        mgr44__std__lane13_strm0_data_valid  ,

            // manager 44, lane 13, stream 1      
            input   wire                                        std__mgr44__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane13_strm1_data        ,
            output  wire                                        mgr44__std__lane13_strm1_data_valid  ,

            // manager 44, lane 14, stream 0      
            input   wire                                        std__mgr44__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane14_strm0_data        ,
            output  wire                                        mgr44__std__lane14_strm0_data_valid  ,

            // manager 44, lane 14, stream 1      
            input   wire                                        std__mgr44__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane14_strm1_data        ,
            output  wire                                        mgr44__std__lane14_strm1_data_valid  ,

            // manager 44, lane 15, stream 0      
            input   wire                                        std__mgr44__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane15_strm0_data        ,
            output  wire                                        mgr44__std__lane15_strm0_data_valid  ,

            // manager 44, lane 15, stream 1      
            input   wire                                        std__mgr44__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane15_strm1_data        ,
            output  wire                                        mgr44__std__lane15_strm1_data_valid  ,

            // manager 44, lane 16, stream 0      
            input   wire                                        std__mgr44__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane16_strm0_data        ,
            output  wire                                        mgr44__std__lane16_strm0_data_valid  ,

            // manager 44, lane 16, stream 1      
            input   wire                                        std__mgr44__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane16_strm1_data        ,
            output  wire                                        mgr44__std__lane16_strm1_data_valid  ,

            // manager 44, lane 17, stream 0      
            input   wire                                        std__mgr44__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane17_strm0_data        ,
            output  wire                                        mgr44__std__lane17_strm0_data_valid  ,

            // manager 44, lane 17, stream 1      
            input   wire                                        std__mgr44__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane17_strm1_data        ,
            output  wire                                        mgr44__std__lane17_strm1_data_valid  ,

            // manager 44, lane 18, stream 0      
            input   wire                                        std__mgr44__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane18_strm0_data        ,
            output  wire                                        mgr44__std__lane18_strm0_data_valid  ,

            // manager 44, lane 18, stream 1      
            input   wire                                        std__mgr44__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane18_strm1_data        ,
            output  wire                                        mgr44__std__lane18_strm1_data_valid  ,

            // manager 44, lane 19, stream 0      
            input   wire                                        std__mgr44__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane19_strm0_data        ,
            output  wire                                        mgr44__std__lane19_strm0_data_valid  ,

            // manager 44, lane 19, stream 1      
            input   wire                                        std__mgr44__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane19_strm1_data        ,
            output  wire                                        mgr44__std__lane19_strm1_data_valid  ,

            // manager 44, lane 20, stream 0      
            input   wire                                        std__mgr44__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane20_strm0_data        ,
            output  wire                                        mgr44__std__lane20_strm0_data_valid  ,

            // manager 44, lane 20, stream 1      
            input   wire                                        std__mgr44__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane20_strm1_data        ,
            output  wire                                        mgr44__std__lane20_strm1_data_valid  ,

            // manager 44, lane 21, stream 0      
            input   wire                                        std__mgr44__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane21_strm0_data        ,
            output  wire                                        mgr44__std__lane21_strm0_data_valid  ,

            // manager 44, lane 21, stream 1      
            input   wire                                        std__mgr44__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane21_strm1_data        ,
            output  wire                                        mgr44__std__lane21_strm1_data_valid  ,

            // manager 44, lane 22, stream 0      
            input   wire                                        std__mgr44__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane22_strm0_data        ,
            output  wire                                        mgr44__std__lane22_strm0_data_valid  ,

            // manager 44, lane 22, stream 1      
            input   wire                                        std__mgr44__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane22_strm1_data        ,
            output  wire                                        mgr44__std__lane22_strm1_data_valid  ,

            // manager 44, lane 23, stream 0      
            input   wire                                        std__mgr44__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane23_strm0_data        ,
            output  wire                                        mgr44__std__lane23_strm0_data_valid  ,

            // manager 44, lane 23, stream 1      
            input   wire                                        std__mgr44__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane23_strm1_data        ,
            output  wire                                        mgr44__std__lane23_strm1_data_valid  ,

            // manager 44, lane 24, stream 0      
            input   wire                                        std__mgr44__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane24_strm0_data        ,
            output  wire                                        mgr44__std__lane24_strm0_data_valid  ,

            // manager 44, lane 24, stream 1      
            input   wire                                        std__mgr44__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane24_strm1_data        ,
            output  wire                                        mgr44__std__lane24_strm1_data_valid  ,

            // manager 44, lane 25, stream 0      
            input   wire                                        std__mgr44__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane25_strm0_data        ,
            output  wire                                        mgr44__std__lane25_strm0_data_valid  ,

            // manager 44, lane 25, stream 1      
            input   wire                                        std__mgr44__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane25_strm1_data        ,
            output  wire                                        mgr44__std__lane25_strm1_data_valid  ,

            // manager 44, lane 26, stream 0      
            input   wire                                        std__mgr44__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane26_strm0_data        ,
            output  wire                                        mgr44__std__lane26_strm0_data_valid  ,

            // manager 44, lane 26, stream 1      
            input   wire                                        std__mgr44__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane26_strm1_data        ,
            output  wire                                        mgr44__std__lane26_strm1_data_valid  ,

            // manager 44, lane 27, stream 0      
            input   wire                                        std__mgr44__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane27_strm0_data        ,
            output  wire                                        mgr44__std__lane27_strm0_data_valid  ,

            // manager 44, lane 27, stream 1      
            input   wire                                        std__mgr44__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane27_strm1_data        ,
            output  wire                                        mgr44__std__lane27_strm1_data_valid  ,

            // manager 44, lane 28, stream 0      
            input   wire                                        std__mgr44__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane28_strm0_data        ,
            output  wire                                        mgr44__std__lane28_strm0_data_valid  ,

            // manager 44, lane 28, stream 1      
            input   wire                                        std__mgr44__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane28_strm1_data        ,
            output  wire                                        mgr44__std__lane28_strm1_data_valid  ,

            // manager 44, lane 29, stream 0      
            input   wire                                        std__mgr44__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane29_strm0_data        ,
            output  wire                                        mgr44__std__lane29_strm0_data_valid  ,

            // manager 44, lane 29, stream 1      
            input   wire                                        std__mgr44__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane29_strm1_data        ,
            output  wire                                        mgr44__std__lane29_strm1_data_valid  ,

            // manager 44, lane 30, stream 0      
            input   wire                                        std__mgr44__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane30_strm0_data        ,
            output  wire                                        mgr44__std__lane30_strm0_data_valid  ,

            // manager 44, lane 30, stream 1      
            input   wire                                        std__mgr44__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane30_strm1_data        ,
            output  wire                                        mgr44__std__lane30_strm1_data_valid  ,

            // manager 44, lane 31, stream 0      
            input   wire                                        std__mgr44__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane31_strm0_data        ,
            output  wire                                        mgr44__std__lane31_strm0_data_valid  ,

            // manager 44, lane 31, stream 1      
            input   wire                                        std__mgr44__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr44__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr44__std__lane31_strm1_data        ,
            output  wire                                        mgr44__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 45, lane 0, stream 0      
            input   wire                                        std__mgr45__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane0_strm0_data        ,
            output  wire                                        mgr45__std__lane0_strm0_data_valid  ,

            // manager 45, lane 0, stream 1      
            input   wire                                        std__mgr45__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane0_strm1_data        ,
            output  wire                                        mgr45__std__lane0_strm1_data_valid  ,

            // manager 45, lane 1, stream 0      
            input   wire                                        std__mgr45__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane1_strm0_data        ,
            output  wire                                        mgr45__std__lane1_strm0_data_valid  ,

            // manager 45, lane 1, stream 1      
            input   wire                                        std__mgr45__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane1_strm1_data        ,
            output  wire                                        mgr45__std__lane1_strm1_data_valid  ,

            // manager 45, lane 2, stream 0      
            input   wire                                        std__mgr45__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane2_strm0_data        ,
            output  wire                                        mgr45__std__lane2_strm0_data_valid  ,

            // manager 45, lane 2, stream 1      
            input   wire                                        std__mgr45__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane2_strm1_data        ,
            output  wire                                        mgr45__std__lane2_strm1_data_valid  ,

            // manager 45, lane 3, stream 0      
            input   wire                                        std__mgr45__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane3_strm0_data        ,
            output  wire                                        mgr45__std__lane3_strm0_data_valid  ,

            // manager 45, lane 3, stream 1      
            input   wire                                        std__mgr45__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane3_strm1_data        ,
            output  wire                                        mgr45__std__lane3_strm1_data_valid  ,

            // manager 45, lane 4, stream 0      
            input   wire                                        std__mgr45__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane4_strm0_data        ,
            output  wire                                        mgr45__std__lane4_strm0_data_valid  ,

            // manager 45, lane 4, stream 1      
            input   wire                                        std__mgr45__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane4_strm1_data        ,
            output  wire                                        mgr45__std__lane4_strm1_data_valid  ,

            // manager 45, lane 5, stream 0      
            input   wire                                        std__mgr45__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane5_strm0_data        ,
            output  wire                                        mgr45__std__lane5_strm0_data_valid  ,

            // manager 45, lane 5, stream 1      
            input   wire                                        std__mgr45__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane5_strm1_data        ,
            output  wire                                        mgr45__std__lane5_strm1_data_valid  ,

            // manager 45, lane 6, stream 0      
            input   wire                                        std__mgr45__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane6_strm0_data        ,
            output  wire                                        mgr45__std__lane6_strm0_data_valid  ,

            // manager 45, lane 6, stream 1      
            input   wire                                        std__mgr45__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane6_strm1_data        ,
            output  wire                                        mgr45__std__lane6_strm1_data_valid  ,

            // manager 45, lane 7, stream 0      
            input   wire                                        std__mgr45__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane7_strm0_data        ,
            output  wire                                        mgr45__std__lane7_strm0_data_valid  ,

            // manager 45, lane 7, stream 1      
            input   wire                                        std__mgr45__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane7_strm1_data        ,
            output  wire                                        mgr45__std__lane7_strm1_data_valid  ,

            // manager 45, lane 8, stream 0      
            input   wire                                        std__mgr45__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane8_strm0_data        ,
            output  wire                                        mgr45__std__lane8_strm0_data_valid  ,

            // manager 45, lane 8, stream 1      
            input   wire                                        std__mgr45__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane8_strm1_data        ,
            output  wire                                        mgr45__std__lane8_strm1_data_valid  ,

            // manager 45, lane 9, stream 0      
            input   wire                                        std__mgr45__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane9_strm0_data        ,
            output  wire                                        mgr45__std__lane9_strm0_data_valid  ,

            // manager 45, lane 9, stream 1      
            input   wire                                        std__mgr45__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane9_strm1_data        ,
            output  wire                                        mgr45__std__lane9_strm1_data_valid  ,

            // manager 45, lane 10, stream 0      
            input   wire                                        std__mgr45__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane10_strm0_data        ,
            output  wire                                        mgr45__std__lane10_strm0_data_valid  ,

            // manager 45, lane 10, stream 1      
            input   wire                                        std__mgr45__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane10_strm1_data        ,
            output  wire                                        mgr45__std__lane10_strm1_data_valid  ,

            // manager 45, lane 11, stream 0      
            input   wire                                        std__mgr45__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane11_strm0_data        ,
            output  wire                                        mgr45__std__lane11_strm0_data_valid  ,

            // manager 45, lane 11, stream 1      
            input   wire                                        std__mgr45__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane11_strm1_data        ,
            output  wire                                        mgr45__std__lane11_strm1_data_valid  ,

            // manager 45, lane 12, stream 0      
            input   wire                                        std__mgr45__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane12_strm0_data        ,
            output  wire                                        mgr45__std__lane12_strm0_data_valid  ,

            // manager 45, lane 12, stream 1      
            input   wire                                        std__mgr45__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane12_strm1_data        ,
            output  wire                                        mgr45__std__lane12_strm1_data_valid  ,

            // manager 45, lane 13, stream 0      
            input   wire                                        std__mgr45__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane13_strm0_data        ,
            output  wire                                        mgr45__std__lane13_strm0_data_valid  ,

            // manager 45, lane 13, stream 1      
            input   wire                                        std__mgr45__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane13_strm1_data        ,
            output  wire                                        mgr45__std__lane13_strm1_data_valid  ,

            // manager 45, lane 14, stream 0      
            input   wire                                        std__mgr45__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane14_strm0_data        ,
            output  wire                                        mgr45__std__lane14_strm0_data_valid  ,

            // manager 45, lane 14, stream 1      
            input   wire                                        std__mgr45__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane14_strm1_data        ,
            output  wire                                        mgr45__std__lane14_strm1_data_valid  ,

            // manager 45, lane 15, stream 0      
            input   wire                                        std__mgr45__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane15_strm0_data        ,
            output  wire                                        mgr45__std__lane15_strm0_data_valid  ,

            // manager 45, lane 15, stream 1      
            input   wire                                        std__mgr45__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane15_strm1_data        ,
            output  wire                                        mgr45__std__lane15_strm1_data_valid  ,

            // manager 45, lane 16, stream 0      
            input   wire                                        std__mgr45__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane16_strm0_data        ,
            output  wire                                        mgr45__std__lane16_strm0_data_valid  ,

            // manager 45, lane 16, stream 1      
            input   wire                                        std__mgr45__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane16_strm1_data        ,
            output  wire                                        mgr45__std__lane16_strm1_data_valid  ,

            // manager 45, lane 17, stream 0      
            input   wire                                        std__mgr45__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane17_strm0_data        ,
            output  wire                                        mgr45__std__lane17_strm0_data_valid  ,

            // manager 45, lane 17, stream 1      
            input   wire                                        std__mgr45__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane17_strm1_data        ,
            output  wire                                        mgr45__std__lane17_strm1_data_valid  ,

            // manager 45, lane 18, stream 0      
            input   wire                                        std__mgr45__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane18_strm0_data        ,
            output  wire                                        mgr45__std__lane18_strm0_data_valid  ,

            // manager 45, lane 18, stream 1      
            input   wire                                        std__mgr45__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane18_strm1_data        ,
            output  wire                                        mgr45__std__lane18_strm1_data_valid  ,

            // manager 45, lane 19, stream 0      
            input   wire                                        std__mgr45__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane19_strm0_data        ,
            output  wire                                        mgr45__std__lane19_strm0_data_valid  ,

            // manager 45, lane 19, stream 1      
            input   wire                                        std__mgr45__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane19_strm1_data        ,
            output  wire                                        mgr45__std__lane19_strm1_data_valid  ,

            // manager 45, lane 20, stream 0      
            input   wire                                        std__mgr45__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane20_strm0_data        ,
            output  wire                                        mgr45__std__lane20_strm0_data_valid  ,

            // manager 45, lane 20, stream 1      
            input   wire                                        std__mgr45__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane20_strm1_data        ,
            output  wire                                        mgr45__std__lane20_strm1_data_valid  ,

            // manager 45, lane 21, stream 0      
            input   wire                                        std__mgr45__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane21_strm0_data        ,
            output  wire                                        mgr45__std__lane21_strm0_data_valid  ,

            // manager 45, lane 21, stream 1      
            input   wire                                        std__mgr45__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane21_strm1_data        ,
            output  wire                                        mgr45__std__lane21_strm1_data_valid  ,

            // manager 45, lane 22, stream 0      
            input   wire                                        std__mgr45__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane22_strm0_data        ,
            output  wire                                        mgr45__std__lane22_strm0_data_valid  ,

            // manager 45, lane 22, stream 1      
            input   wire                                        std__mgr45__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane22_strm1_data        ,
            output  wire                                        mgr45__std__lane22_strm1_data_valid  ,

            // manager 45, lane 23, stream 0      
            input   wire                                        std__mgr45__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane23_strm0_data        ,
            output  wire                                        mgr45__std__lane23_strm0_data_valid  ,

            // manager 45, lane 23, stream 1      
            input   wire                                        std__mgr45__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane23_strm1_data        ,
            output  wire                                        mgr45__std__lane23_strm1_data_valid  ,

            // manager 45, lane 24, stream 0      
            input   wire                                        std__mgr45__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane24_strm0_data        ,
            output  wire                                        mgr45__std__lane24_strm0_data_valid  ,

            // manager 45, lane 24, stream 1      
            input   wire                                        std__mgr45__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane24_strm1_data        ,
            output  wire                                        mgr45__std__lane24_strm1_data_valid  ,

            // manager 45, lane 25, stream 0      
            input   wire                                        std__mgr45__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane25_strm0_data        ,
            output  wire                                        mgr45__std__lane25_strm0_data_valid  ,

            // manager 45, lane 25, stream 1      
            input   wire                                        std__mgr45__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane25_strm1_data        ,
            output  wire                                        mgr45__std__lane25_strm1_data_valid  ,

            // manager 45, lane 26, stream 0      
            input   wire                                        std__mgr45__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane26_strm0_data        ,
            output  wire                                        mgr45__std__lane26_strm0_data_valid  ,

            // manager 45, lane 26, stream 1      
            input   wire                                        std__mgr45__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane26_strm1_data        ,
            output  wire                                        mgr45__std__lane26_strm1_data_valid  ,

            // manager 45, lane 27, stream 0      
            input   wire                                        std__mgr45__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane27_strm0_data        ,
            output  wire                                        mgr45__std__lane27_strm0_data_valid  ,

            // manager 45, lane 27, stream 1      
            input   wire                                        std__mgr45__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane27_strm1_data        ,
            output  wire                                        mgr45__std__lane27_strm1_data_valid  ,

            // manager 45, lane 28, stream 0      
            input   wire                                        std__mgr45__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane28_strm0_data        ,
            output  wire                                        mgr45__std__lane28_strm0_data_valid  ,

            // manager 45, lane 28, stream 1      
            input   wire                                        std__mgr45__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane28_strm1_data        ,
            output  wire                                        mgr45__std__lane28_strm1_data_valid  ,

            // manager 45, lane 29, stream 0      
            input   wire                                        std__mgr45__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane29_strm0_data        ,
            output  wire                                        mgr45__std__lane29_strm0_data_valid  ,

            // manager 45, lane 29, stream 1      
            input   wire                                        std__mgr45__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane29_strm1_data        ,
            output  wire                                        mgr45__std__lane29_strm1_data_valid  ,

            // manager 45, lane 30, stream 0      
            input   wire                                        std__mgr45__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane30_strm0_data        ,
            output  wire                                        mgr45__std__lane30_strm0_data_valid  ,

            // manager 45, lane 30, stream 1      
            input   wire                                        std__mgr45__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane30_strm1_data        ,
            output  wire                                        mgr45__std__lane30_strm1_data_valid  ,

            // manager 45, lane 31, stream 0      
            input   wire                                        std__mgr45__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane31_strm0_data        ,
            output  wire                                        mgr45__std__lane31_strm0_data_valid  ,

            // manager 45, lane 31, stream 1      
            input   wire                                        std__mgr45__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr45__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr45__std__lane31_strm1_data        ,
            output  wire                                        mgr45__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 46, lane 0, stream 0      
            input   wire                                        std__mgr46__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane0_strm0_data        ,
            output  wire                                        mgr46__std__lane0_strm0_data_valid  ,

            // manager 46, lane 0, stream 1      
            input   wire                                        std__mgr46__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane0_strm1_data        ,
            output  wire                                        mgr46__std__lane0_strm1_data_valid  ,

            // manager 46, lane 1, stream 0      
            input   wire                                        std__mgr46__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane1_strm0_data        ,
            output  wire                                        mgr46__std__lane1_strm0_data_valid  ,

            // manager 46, lane 1, stream 1      
            input   wire                                        std__mgr46__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane1_strm1_data        ,
            output  wire                                        mgr46__std__lane1_strm1_data_valid  ,

            // manager 46, lane 2, stream 0      
            input   wire                                        std__mgr46__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane2_strm0_data        ,
            output  wire                                        mgr46__std__lane2_strm0_data_valid  ,

            // manager 46, lane 2, stream 1      
            input   wire                                        std__mgr46__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane2_strm1_data        ,
            output  wire                                        mgr46__std__lane2_strm1_data_valid  ,

            // manager 46, lane 3, stream 0      
            input   wire                                        std__mgr46__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane3_strm0_data        ,
            output  wire                                        mgr46__std__lane3_strm0_data_valid  ,

            // manager 46, lane 3, stream 1      
            input   wire                                        std__mgr46__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane3_strm1_data        ,
            output  wire                                        mgr46__std__lane3_strm1_data_valid  ,

            // manager 46, lane 4, stream 0      
            input   wire                                        std__mgr46__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane4_strm0_data        ,
            output  wire                                        mgr46__std__lane4_strm0_data_valid  ,

            // manager 46, lane 4, stream 1      
            input   wire                                        std__mgr46__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane4_strm1_data        ,
            output  wire                                        mgr46__std__lane4_strm1_data_valid  ,

            // manager 46, lane 5, stream 0      
            input   wire                                        std__mgr46__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane5_strm0_data        ,
            output  wire                                        mgr46__std__lane5_strm0_data_valid  ,

            // manager 46, lane 5, stream 1      
            input   wire                                        std__mgr46__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane5_strm1_data        ,
            output  wire                                        mgr46__std__lane5_strm1_data_valid  ,

            // manager 46, lane 6, stream 0      
            input   wire                                        std__mgr46__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane6_strm0_data        ,
            output  wire                                        mgr46__std__lane6_strm0_data_valid  ,

            // manager 46, lane 6, stream 1      
            input   wire                                        std__mgr46__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane6_strm1_data        ,
            output  wire                                        mgr46__std__lane6_strm1_data_valid  ,

            // manager 46, lane 7, stream 0      
            input   wire                                        std__mgr46__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane7_strm0_data        ,
            output  wire                                        mgr46__std__lane7_strm0_data_valid  ,

            // manager 46, lane 7, stream 1      
            input   wire                                        std__mgr46__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane7_strm1_data        ,
            output  wire                                        mgr46__std__lane7_strm1_data_valid  ,

            // manager 46, lane 8, stream 0      
            input   wire                                        std__mgr46__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane8_strm0_data        ,
            output  wire                                        mgr46__std__lane8_strm0_data_valid  ,

            // manager 46, lane 8, stream 1      
            input   wire                                        std__mgr46__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane8_strm1_data        ,
            output  wire                                        mgr46__std__lane8_strm1_data_valid  ,

            // manager 46, lane 9, stream 0      
            input   wire                                        std__mgr46__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane9_strm0_data        ,
            output  wire                                        mgr46__std__lane9_strm0_data_valid  ,

            // manager 46, lane 9, stream 1      
            input   wire                                        std__mgr46__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane9_strm1_data        ,
            output  wire                                        mgr46__std__lane9_strm1_data_valid  ,

            // manager 46, lane 10, stream 0      
            input   wire                                        std__mgr46__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane10_strm0_data        ,
            output  wire                                        mgr46__std__lane10_strm0_data_valid  ,

            // manager 46, lane 10, stream 1      
            input   wire                                        std__mgr46__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane10_strm1_data        ,
            output  wire                                        mgr46__std__lane10_strm1_data_valid  ,

            // manager 46, lane 11, stream 0      
            input   wire                                        std__mgr46__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane11_strm0_data        ,
            output  wire                                        mgr46__std__lane11_strm0_data_valid  ,

            // manager 46, lane 11, stream 1      
            input   wire                                        std__mgr46__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane11_strm1_data        ,
            output  wire                                        mgr46__std__lane11_strm1_data_valid  ,

            // manager 46, lane 12, stream 0      
            input   wire                                        std__mgr46__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane12_strm0_data        ,
            output  wire                                        mgr46__std__lane12_strm0_data_valid  ,

            // manager 46, lane 12, stream 1      
            input   wire                                        std__mgr46__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane12_strm1_data        ,
            output  wire                                        mgr46__std__lane12_strm1_data_valid  ,

            // manager 46, lane 13, stream 0      
            input   wire                                        std__mgr46__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane13_strm0_data        ,
            output  wire                                        mgr46__std__lane13_strm0_data_valid  ,

            // manager 46, lane 13, stream 1      
            input   wire                                        std__mgr46__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane13_strm1_data        ,
            output  wire                                        mgr46__std__lane13_strm1_data_valid  ,

            // manager 46, lane 14, stream 0      
            input   wire                                        std__mgr46__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane14_strm0_data        ,
            output  wire                                        mgr46__std__lane14_strm0_data_valid  ,

            // manager 46, lane 14, stream 1      
            input   wire                                        std__mgr46__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane14_strm1_data        ,
            output  wire                                        mgr46__std__lane14_strm1_data_valid  ,

            // manager 46, lane 15, stream 0      
            input   wire                                        std__mgr46__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane15_strm0_data        ,
            output  wire                                        mgr46__std__lane15_strm0_data_valid  ,

            // manager 46, lane 15, stream 1      
            input   wire                                        std__mgr46__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane15_strm1_data        ,
            output  wire                                        mgr46__std__lane15_strm1_data_valid  ,

            // manager 46, lane 16, stream 0      
            input   wire                                        std__mgr46__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane16_strm0_data        ,
            output  wire                                        mgr46__std__lane16_strm0_data_valid  ,

            // manager 46, lane 16, stream 1      
            input   wire                                        std__mgr46__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane16_strm1_data        ,
            output  wire                                        mgr46__std__lane16_strm1_data_valid  ,

            // manager 46, lane 17, stream 0      
            input   wire                                        std__mgr46__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane17_strm0_data        ,
            output  wire                                        mgr46__std__lane17_strm0_data_valid  ,

            // manager 46, lane 17, stream 1      
            input   wire                                        std__mgr46__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane17_strm1_data        ,
            output  wire                                        mgr46__std__lane17_strm1_data_valid  ,

            // manager 46, lane 18, stream 0      
            input   wire                                        std__mgr46__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane18_strm0_data        ,
            output  wire                                        mgr46__std__lane18_strm0_data_valid  ,

            // manager 46, lane 18, stream 1      
            input   wire                                        std__mgr46__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane18_strm1_data        ,
            output  wire                                        mgr46__std__lane18_strm1_data_valid  ,

            // manager 46, lane 19, stream 0      
            input   wire                                        std__mgr46__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane19_strm0_data        ,
            output  wire                                        mgr46__std__lane19_strm0_data_valid  ,

            // manager 46, lane 19, stream 1      
            input   wire                                        std__mgr46__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane19_strm1_data        ,
            output  wire                                        mgr46__std__lane19_strm1_data_valid  ,

            // manager 46, lane 20, stream 0      
            input   wire                                        std__mgr46__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane20_strm0_data        ,
            output  wire                                        mgr46__std__lane20_strm0_data_valid  ,

            // manager 46, lane 20, stream 1      
            input   wire                                        std__mgr46__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane20_strm1_data        ,
            output  wire                                        mgr46__std__lane20_strm1_data_valid  ,

            // manager 46, lane 21, stream 0      
            input   wire                                        std__mgr46__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane21_strm0_data        ,
            output  wire                                        mgr46__std__lane21_strm0_data_valid  ,

            // manager 46, lane 21, stream 1      
            input   wire                                        std__mgr46__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane21_strm1_data        ,
            output  wire                                        mgr46__std__lane21_strm1_data_valid  ,

            // manager 46, lane 22, stream 0      
            input   wire                                        std__mgr46__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane22_strm0_data        ,
            output  wire                                        mgr46__std__lane22_strm0_data_valid  ,

            // manager 46, lane 22, stream 1      
            input   wire                                        std__mgr46__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane22_strm1_data        ,
            output  wire                                        mgr46__std__lane22_strm1_data_valid  ,

            // manager 46, lane 23, stream 0      
            input   wire                                        std__mgr46__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane23_strm0_data        ,
            output  wire                                        mgr46__std__lane23_strm0_data_valid  ,

            // manager 46, lane 23, stream 1      
            input   wire                                        std__mgr46__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane23_strm1_data        ,
            output  wire                                        mgr46__std__lane23_strm1_data_valid  ,

            // manager 46, lane 24, stream 0      
            input   wire                                        std__mgr46__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane24_strm0_data        ,
            output  wire                                        mgr46__std__lane24_strm0_data_valid  ,

            // manager 46, lane 24, stream 1      
            input   wire                                        std__mgr46__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane24_strm1_data        ,
            output  wire                                        mgr46__std__lane24_strm1_data_valid  ,

            // manager 46, lane 25, stream 0      
            input   wire                                        std__mgr46__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane25_strm0_data        ,
            output  wire                                        mgr46__std__lane25_strm0_data_valid  ,

            // manager 46, lane 25, stream 1      
            input   wire                                        std__mgr46__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane25_strm1_data        ,
            output  wire                                        mgr46__std__lane25_strm1_data_valid  ,

            // manager 46, lane 26, stream 0      
            input   wire                                        std__mgr46__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane26_strm0_data        ,
            output  wire                                        mgr46__std__lane26_strm0_data_valid  ,

            // manager 46, lane 26, stream 1      
            input   wire                                        std__mgr46__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane26_strm1_data        ,
            output  wire                                        mgr46__std__lane26_strm1_data_valid  ,

            // manager 46, lane 27, stream 0      
            input   wire                                        std__mgr46__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane27_strm0_data        ,
            output  wire                                        mgr46__std__lane27_strm0_data_valid  ,

            // manager 46, lane 27, stream 1      
            input   wire                                        std__mgr46__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane27_strm1_data        ,
            output  wire                                        mgr46__std__lane27_strm1_data_valid  ,

            // manager 46, lane 28, stream 0      
            input   wire                                        std__mgr46__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane28_strm0_data        ,
            output  wire                                        mgr46__std__lane28_strm0_data_valid  ,

            // manager 46, lane 28, stream 1      
            input   wire                                        std__mgr46__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane28_strm1_data        ,
            output  wire                                        mgr46__std__lane28_strm1_data_valid  ,

            // manager 46, lane 29, stream 0      
            input   wire                                        std__mgr46__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane29_strm0_data        ,
            output  wire                                        mgr46__std__lane29_strm0_data_valid  ,

            // manager 46, lane 29, stream 1      
            input   wire                                        std__mgr46__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane29_strm1_data        ,
            output  wire                                        mgr46__std__lane29_strm1_data_valid  ,

            // manager 46, lane 30, stream 0      
            input   wire                                        std__mgr46__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane30_strm0_data        ,
            output  wire                                        mgr46__std__lane30_strm0_data_valid  ,

            // manager 46, lane 30, stream 1      
            input   wire                                        std__mgr46__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane30_strm1_data        ,
            output  wire                                        mgr46__std__lane30_strm1_data_valid  ,

            // manager 46, lane 31, stream 0      
            input   wire                                        std__mgr46__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane31_strm0_data        ,
            output  wire                                        mgr46__std__lane31_strm0_data_valid  ,

            // manager 46, lane 31, stream 1      
            input   wire                                        std__mgr46__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr46__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr46__std__lane31_strm1_data        ,
            output  wire                                        mgr46__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 47, lane 0, stream 0      
            input   wire                                        std__mgr47__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane0_strm0_data        ,
            output  wire                                        mgr47__std__lane0_strm0_data_valid  ,

            // manager 47, lane 0, stream 1      
            input   wire                                        std__mgr47__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane0_strm1_data        ,
            output  wire                                        mgr47__std__lane0_strm1_data_valid  ,

            // manager 47, lane 1, stream 0      
            input   wire                                        std__mgr47__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane1_strm0_data        ,
            output  wire                                        mgr47__std__lane1_strm0_data_valid  ,

            // manager 47, lane 1, stream 1      
            input   wire                                        std__mgr47__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane1_strm1_data        ,
            output  wire                                        mgr47__std__lane1_strm1_data_valid  ,

            // manager 47, lane 2, stream 0      
            input   wire                                        std__mgr47__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane2_strm0_data        ,
            output  wire                                        mgr47__std__lane2_strm0_data_valid  ,

            // manager 47, lane 2, stream 1      
            input   wire                                        std__mgr47__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane2_strm1_data        ,
            output  wire                                        mgr47__std__lane2_strm1_data_valid  ,

            // manager 47, lane 3, stream 0      
            input   wire                                        std__mgr47__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane3_strm0_data        ,
            output  wire                                        mgr47__std__lane3_strm0_data_valid  ,

            // manager 47, lane 3, stream 1      
            input   wire                                        std__mgr47__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane3_strm1_data        ,
            output  wire                                        mgr47__std__lane3_strm1_data_valid  ,

            // manager 47, lane 4, stream 0      
            input   wire                                        std__mgr47__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane4_strm0_data        ,
            output  wire                                        mgr47__std__lane4_strm0_data_valid  ,

            // manager 47, lane 4, stream 1      
            input   wire                                        std__mgr47__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane4_strm1_data        ,
            output  wire                                        mgr47__std__lane4_strm1_data_valid  ,

            // manager 47, lane 5, stream 0      
            input   wire                                        std__mgr47__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane5_strm0_data        ,
            output  wire                                        mgr47__std__lane5_strm0_data_valid  ,

            // manager 47, lane 5, stream 1      
            input   wire                                        std__mgr47__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane5_strm1_data        ,
            output  wire                                        mgr47__std__lane5_strm1_data_valid  ,

            // manager 47, lane 6, stream 0      
            input   wire                                        std__mgr47__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane6_strm0_data        ,
            output  wire                                        mgr47__std__lane6_strm0_data_valid  ,

            // manager 47, lane 6, stream 1      
            input   wire                                        std__mgr47__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane6_strm1_data        ,
            output  wire                                        mgr47__std__lane6_strm1_data_valid  ,

            // manager 47, lane 7, stream 0      
            input   wire                                        std__mgr47__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane7_strm0_data        ,
            output  wire                                        mgr47__std__lane7_strm0_data_valid  ,

            // manager 47, lane 7, stream 1      
            input   wire                                        std__mgr47__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane7_strm1_data        ,
            output  wire                                        mgr47__std__lane7_strm1_data_valid  ,

            // manager 47, lane 8, stream 0      
            input   wire                                        std__mgr47__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane8_strm0_data        ,
            output  wire                                        mgr47__std__lane8_strm0_data_valid  ,

            // manager 47, lane 8, stream 1      
            input   wire                                        std__mgr47__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane8_strm1_data        ,
            output  wire                                        mgr47__std__lane8_strm1_data_valid  ,

            // manager 47, lane 9, stream 0      
            input   wire                                        std__mgr47__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane9_strm0_data        ,
            output  wire                                        mgr47__std__lane9_strm0_data_valid  ,

            // manager 47, lane 9, stream 1      
            input   wire                                        std__mgr47__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane9_strm1_data        ,
            output  wire                                        mgr47__std__lane9_strm1_data_valid  ,

            // manager 47, lane 10, stream 0      
            input   wire                                        std__mgr47__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane10_strm0_data        ,
            output  wire                                        mgr47__std__lane10_strm0_data_valid  ,

            // manager 47, lane 10, stream 1      
            input   wire                                        std__mgr47__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane10_strm1_data        ,
            output  wire                                        mgr47__std__lane10_strm1_data_valid  ,

            // manager 47, lane 11, stream 0      
            input   wire                                        std__mgr47__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane11_strm0_data        ,
            output  wire                                        mgr47__std__lane11_strm0_data_valid  ,

            // manager 47, lane 11, stream 1      
            input   wire                                        std__mgr47__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane11_strm1_data        ,
            output  wire                                        mgr47__std__lane11_strm1_data_valid  ,

            // manager 47, lane 12, stream 0      
            input   wire                                        std__mgr47__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane12_strm0_data        ,
            output  wire                                        mgr47__std__lane12_strm0_data_valid  ,

            // manager 47, lane 12, stream 1      
            input   wire                                        std__mgr47__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane12_strm1_data        ,
            output  wire                                        mgr47__std__lane12_strm1_data_valid  ,

            // manager 47, lane 13, stream 0      
            input   wire                                        std__mgr47__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane13_strm0_data        ,
            output  wire                                        mgr47__std__lane13_strm0_data_valid  ,

            // manager 47, lane 13, stream 1      
            input   wire                                        std__mgr47__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane13_strm1_data        ,
            output  wire                                        mgr47__std__lane13_strm1_data_valid  ,

            // manager 47, lane 14, stream 0      
            input   wire                                        std__mgr47__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane14_strm0_data        ,
            output  wire                                        mgr47__std__lane14_strm0_data_valid  ,

            // manager 47, lane 14, stream 1      
            input   wire                                        std__mgr47__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane14_strm1_data        ,
            output  wire                                        mgr47__std__lane14_strm1_data_valid  ,

            // manager 47, lane 15, stream 0      
            input   wire                                        std__mgr47__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane15_strm0_data        ,
            output  wire                                        mgr47__std__lane15_strm0_data_valid  ,

            // manager 47, lane 15, stream 1      
            input   wire                                        std__mgr47__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane15_strm1_data        ,
            output  wire                                        mgr47__std__lane15_strm1_data_valid  ,

            // manager 47, lane 16, stream 0      
            input   wire                                        std__mgr47__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane16_strm0_data        ,
            output  wire                                        mgr47__std__lane16_strm0_data_valid  ,

            // manager 47, lane 16, stream 1      
            input   wire                                        std__mgr47__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane16_strm1_data        ,
            output  wire                                        mgr47__std__lane16_strm1_data_valid  ,

            // manager 47, lane 17, stream 0      
            input   wire                                        std__mgr47__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane17_strm0_data        ,
            output  wire                                        mgr47__std__lane17_strm0_data_valid  ,

            // manager 47, lane 17, stream 1      
            input   wire                                        std__mgr47__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane17_strm1_data        ,
            output  wire                                        mgr47__std__lane17_strm1_data_valid  ,

            // manager 47, lane 18, stream 0      
            input   wire                                        std__mgr47__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane18_strm0_data        ,
            output  wire                                        mgr47__std__lane18_strm0_data_valid  ,

            // manager 47, lane 18, stream 1      
            input   wire                                        std__mgr47__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane18_strm1_data        ,
            output  wire                                        mgr47__std__lane18_strm1_data_valid  ,

            // manager 47, lane 19, stream 0      
            input   wire                                        std__mgr47__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane19_strm0_data        ,
            output  wire                                        mgr47__std__lane19_strm0_data_valid  ,

            // manager 47, lane 19, stream 1      
            input   wire                                        std__mgr47__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane19_strm1_data        ,
            output  wire                                        mgr47__std__lane19_strm1_data_valid  ,

            // manager 47, lane 20, stream 0      
            input   wire                                        std__mgr47__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane20_strm0_data        ,
            output  wire                                        mgr47__std__lane20_strm0_data_valid  ,

            // manager 47, lane 20, stream 1      
            input   wire                                        std__mgr47__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane20_strm1_data        ,
            output  wire                                        mgr47__std__lane20_strm1_data_valid  ,

            // manager 47, lane 21, stream 0      
            input   wire                                        std__mgr47__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane21_strm0_data        ,
            output  wire                                        mgr47__std__lane21_strm0_data_valid  ,

            // manager 47, lane 21, stream 1      
            input   wire                                        std__mgr47__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane21_strm1_data        ,
            output  wire                                        mgr47__std__lane21_strm1_data_valid  ,

            // manager 47, lane 22, stream 0      
            input   wire                                        std__mgr47__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane22_strm0_data        ,
            output  wire                                        mgr47__std__lane22_strm0_data_valid  ,

            // manager 47, lane 22, stream 1      
            input   wire                                        std__mgr47__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane22_strm1_data        ,
            output  wire                                        mgr47__std__lane22_strm1_data_valid  ,

            // manager 47, lane 23, stream 0      
            input   wire                                        std__mgr47__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane23_strm0_data        ,
            output  wire                                        mgr47__std__lane23_strm0_data_valid  ,

            // manager 47, lane 23, stream 1      
            input   wire                                        std__mgr47__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane23_strm1_data        ,
            output  wire                                        mgr47__std__lane23_strm1_data_valid  ,

            // manager 47, lane 24, stream 0      
            input   wire                                        std__mgr47__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane24_strm0_data        ,
            output  wire                                        mgr47__std__lane24_strm0_data_valid  ,

            // manager 47, lane 24, stream 1      
            input   wire                                        std__mgr47__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane24_strm1_data        ,
            output  wire                                        mgr47__std__lane24_strm1_data_valid  ,

            // manager 47, lane 25, stream 0      
            input   wire                                        std__mgr47__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane25_strm0_data        ,
            output  wire                                        mgr47__std__lane25_strm0_data_valid  ,

            // manager 47, lane 25, stream 1      
            input   wire                                        std__mgr47__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane25_strm1_data        ,
            output  wire                                        mgr47__std__lane25_strm1_data_valid  ,

            // manager 47, lane 26, stream 0      
            input   wire                                        std__mgr47__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane26_strm0_data        ,
            output  wire                                        mgr47__std__lane26_strm0_data_valid  ,

            // manager 47, lane 26, stream 1      
            input   wire                                        std__mgr47__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane26_strm1_data        ,
            output  wire                                        mgr47__std__lane26_strm1_data_valid  ,

            // manager 47, lane 27, stream 0      
            input   wire                                        std__mgr47__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane27_strm0_data        ,
            output  wire                                        mgr47__std__lane27_strm0_data_valid  ,

            // manager 47, lane 27, stream 1      
            input   wire                                        std__mgr47__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane27_strm1_data        ,
            output  wire                                        mgr47__std__lane27_strm1_data_valid  ,

            // manager 47, lane 28, stream 0      
            input   wire                                        std__mgr47__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane28_strm0_data        ,
            output  wire                                        mgr47__std__lane28_strm0_data_valid  ,

            // manager 47, lane 28, stream 1      
            input   wire                                        std__mgr47__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane28_strm1_data        ,
            output  wire                                        mgr47__std__lane28_strm1_data_valid  ,

            // manager 47, lane 29, stream 0      
            input   wire                                        std__mgr47__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane29_strm0_data        ,
            output  wire                                        mgr47__std__lane29_strm0_data_valid  ,

            // manager 47, lane 29, stream 1      
            input   wire                                        std__mgr47__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane29_strm1_data        ,
            output  wire                                        mgr47__std__lane29_strm1_data_valid  ,

            // manager 47, lane 30, stream 0      
            input   wire                                        std__mgr47__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane30_strm0_data        ,
            output  wire                                        mgr47__std__lane30_strm0_data_valid  ,

            // manager 47, lane 30, stream 1      
            input   wire                                        std__mgr47__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane30_strm1_data        ,
            output  wire                                        mgr47__std__lane30_strm1_data_valid  ,

            // manager 47, lane 31, stream 0      
            input   wire                                        std__mgr47__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane31_strm0_data        ,
            output  wire                                        mgr47__std__lane31_strm0_data_valid  ,

            // manager 47, lane 31, stream 1      
            input   wire                                        std__mgr47__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr47__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr47__std__lane31_strm1_data        ,
            output  wire                                        mgr47__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 48, lane 0, stream 0      
            input   wire                                        std__mgr48__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane0_strm0_data        ,
            output  wire                                        mgr48__std__lane0_strm0_data_valid  ,

            // manager 48, lane 0, stream 1      
            input   wire                                        std__mgr48__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane0_strm1_data        ,
            output  wire                                        mgr48__std__lane0_strm1_data_valid  ,

            // manager 48, lane 1, stream 0      
            input   wire                                        std__mgr48__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane1_strm0_data        ,
            output  wire                                        mgr48__std__lane1_strm0_data_valid  ,

            // manager 48, lane 1, stream 1      
            input   wire                                        std__mgr48__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane1_strm1_data        ,
            output  wire                                        mgr48__std__lane1_strm1_data_valid  ,

            // manager 48, lane 2, stream 0      
            input   wire                                        std__mgr48__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane2_strm0_data        ,
            output  wire                                        mgr48__std__lane2_strm0_data_valid  ,

            // manager 48, lane 2, stream 1      
            input   wire                                        std__mgr48__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane2_strm1_data        ,
            output  wire                                        mgr48__std__lane2_strm1_data_valid  ,

            // manager 48, lane 3, stream 0      
            input   wire                                        std__mgr48__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane3_strm0_data        ,
            output  wire                                        mgr48__std__lane3_strm0_data_valid  ,

            // manager 48, lane 3, stream 1      
            input   wire                                        std__mgr48__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane3_strm1_data        ,
            output  wire                                        mgr48__std__lane3_strm1_data_valid  ,

            // manager 48, lane 4, stream 0      
            input   wire                                        std__mgr48__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane4_strm0_data        ,
            output  wire                                        mgr48__std__lane4_strm0_data_valid  ,

            // manager 48, lane 4, stream 1      
            input   wire                                        std__mgr48__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane4_strm1_data        ,
            output  wire                                        mgr48__std__lane4_strm1_data_valid  ,

            // manager 48, lane 5, stream 0      
            input   wire                                        std__mgr48__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane5_strm0_data        ,
            output  wire                                        mgr48__std__lane5_strm0_data_valid  ,

            // manager 48, lane 5, stream 1      
            input   wire                                        std__mgr48__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane5_strm1_data        ,
            output  wire                                        mgr48__std__lane5_strm1_data_valid  ,

            // manager 48, lane 6, stream 0      
            input   wire                                        std__mgr48__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane6_strm0_data        ,
            output  wire                                        mgr48__std__lane6_strm0_data_valid  ,

            // manager 48, lane 6, stream 1      
            input   wire                                        std__mgr48__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane6_strm1_data        ,
            output  wire                                        mgr48__std__lane6_strm1_data_valid  ,

            // manager 48, lane 7, stream 0      
            input   wire                                        std__mgr48__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane7_strm0_data        ,
            output  wire                                        mgr48__std__lane7_strm0_data_valid  ,

            // manager 48, lane 7, stream 1      
            input   wire                                        std__mgr48__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane7_strm1_data        ,
            output  wire                                        mgr48__std__lane7_strm1_data_valid  ,

            // manager 48, lane 8, stream 0      
            input   wire                                        std__mgr48__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane8_strm0_data        ,
            output  wire                                        mgr48__std__lane8_strm0_data_valid  ,

            // manager 48, lane 8, stream 1      
            input   wire                                        std__mgr48__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane8_strm1_data        ,
            output  wire                                        mgr48__std__lane8_strm1_data_valid  ,

            // manager 48, lane 9, stream 0      
            input   wire                                        std__mgr48__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane9_strm0_data        ,
            output  wire                                        mgr48__std__lane9_strm0_data_valid  ,

            // manager 48, lane 9, stream 1      
            input   wire                                        std__mgr48__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane9_strm1_data        ,
            output  wire                                        mgr48__std__lane9_strm1_data_valid  ,

            // manager 48, lane 10, stream 0      
            input   wire                                        std__mgr48__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane10_strm0_data        ,
            output  wire                                        mgr48__std__lane10_strm0_data_valid  ,

            // manager 48, lane 10, stream 1      
            input   wire                                        std__mgr48__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane10_strm1_data        ,
            output  wire                                        mgr48__std__lane10_strm1_data_valid  ,

            // manager 48, lane 11, stream 0      
            input   wire                                        std__mgr48__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane11_strm0_data        ,
            output  wire                                        mgr48__std__lane11_strm0_data_valid  ,

            // manager 48, lane 11, stream 1      
            input   wire                                        std__mgr48__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane11_strm1_data        ,
            output  wire                                        mgr48__std__lane11_strm1_data_valid  ,

            // manager 48, lane 12, stream 0      
            input   wire                                        std__mgr48__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane12_strm0_data        ,
            output  wire                                        mgr48__std__lane12_strm0_data_valid  ,

            // manager 48, lane 12, stream 1      
            input   wire                                        std__mgr48__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane12_strm1_data        ,
            output  wire                                        mgr48__std__lane12_strm1_data_valid  ,

            // manager 48, lane 13, stream 0      
            input   wire                                        std__mgr48__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane13_strm0_data        ,
            output  wire                                        mgr48__std__lane13_strm0_data_valid  ,

            // manager 48, lane 13, stream 1      
            input   wire                                        std__mgr48__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane13_strm1_data        ,
            output  wire                                        mgr48__std__lane13_strm1_data_valid  ,

            // manager 48, lane 14, stream 0      
            input   wire                                        std__mgr48__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane14_strm0_data        ,
            output  wire                                        mgr48__std__lane14_strm0_data_valid  ,

            // manager 48, lane 14, stream 1      
            input   wire                                        std__mgr48__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane14_strm1_data        ,
            output  wire                                        mgr48__std__lane14_strm1_data_valid  ,

            // manager 48, lane 15, stream 0      
            input   wire                                        std__mgr48__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane15_strm0_data        ,
            output  wire                                        mgr48__std__lane15_strm0_data_valid  ,

            // manager 48, lane 15, stream 1      
            input   wire                                        std__mgr48__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane15_strm1_data        ,
            output  wire                                        mgr48__std__lane15_strm1_data_valid  ,

            // manager 48, lane 16, stream 0      
            input   wire                                        std__mgr48__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane16_strm0_data        ,
            output  wire                                        mgr48__std__lane16_strm0_data_valid  ,

            // manager 48, lane 16, stream 1      
            input   wire                                        std__mgr48__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane16_strm1_data        ,
            output  wire                                        mgr48__std__lane16_strm1_data_valid  ,

            // manager 48, lane 17, stream 0      
            input   wire                                        std__mgr48__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane17_strm0_data        ,
            output  wire                                        mgr48__std__lane17_strm0_data_valid  ,

            // manager 48, lane 17, stream 1      
            input   wire                                        std__mgr48__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane17_strm1_data        ,
            output  wire                                        mgr48__std__lane17_strm1_data_valid  ,

            // manager 48, lane 18, stream 0      
            input   wire                                        std__mgr48__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane18_strm0_data        ,
            output  wire                                        mgr48__std__lane18_strm0_data_valid  ,

            // manager 48, lane 18, stream 1      
            input   wire                                        std__mgr48__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane18_strm1_data        ,
            output  wire                                        mgr48__std__lane18_strm1_data_valid  ,

            // manager 48, lane 19, stream 0      
            input   wire                                        std__mgr48__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane19_strm0_data        ,
            output  wire                                        mgr48__std__lane19_strm0_data_valid  ,

            // manager 48, lane 19, stream 1      
            input   wire                                        std__mgr48__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane19_strm1_data        ,
            output  wire                                        mgr48__std__lane19_strm1_data_valid  ,

            // manager 48, lane 20, stream 0      
            input   wire                                        std__mgr48__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane20_strm0_data        ,
            output  wire                                        mgr48__std__lane20_strm0_data_valid  ,

            // manager 48, lane 20, stream 1      
            input   wire                                        std__mgr48__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane20_strm1_data        ,
            output  wire                                        mgr48__std__lane20_strm1_data_valid  ,

            // manager 48, lane 21, stream 0      
            input   wire                                        std__mgr48__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane21_strm0_data        ,
            output  wire                                        mgr48__std__lane21_strm0_data_valid  ,

            // manager 48, lane 21, stream 1      
            input   wire                                        std__mgr48__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane21_strm1_data        ,
            output  wire                                        mgr48__std__lane21_strm1_data_valid  ,

            // manager 48, lane 22, stream 0      
            input   wire                                        std__mgr48__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane22_strm0_data        ,
            output  wire                                        mgr48__std__lane22_strm0_data_valid  ,

            // manager 48, lane 22, stream 1      
            input   wire                                        std__mgr48__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane22_strm1_data        ,
            output  wire                                        mgr48__std__lane22_strm1_data_valid  ,

            // manager 48, lane 23, stream 0      
            input   wire                                        std__mgr48__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane23_strm0_data        ,
            output  wire                                        mgr48__std__lane23_strm0_data_valid  ,

            // manager 48, lane 23, stream 1      
            input   wire                                        std__mgr48__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane23_strm1_data        ,
            output  wire                                        mgr48__std__lane23_strm1_data_valid  ,

            // manager 48, lane 24, stream 0      
            input   wire                                        std__mgr48__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane24_strm0_data        ,
            output  wire                                        mgr48__std__lane24_strm0_data_valid  ,

            // manager 48, lane 24, stream 1      
            input   wire                                        std__mgr48__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane24_strm1_data        ,
            output  wire                                        mgr48__std__lane24_strm1_data_valid  ,

            // manager 48, lane 25, stream 0      
            input   wire                                        std__mgr48__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane25_strm0_data        ,
            output  wire                                        mgr48__std__lane25_strm0_data_valid  ,

            // manager 48, lane 25, stream 1      
            input   wire                                        std__mgr48__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane25_strm1_data        ,
            output  wire                                        mgr48__std__lane25_strm1_data_valid  ,

            // manager 48, lane 26, stream 0      
            input   wire                                        std__mgr48__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane26_strm0_data        ,
            output  wire                                        mgr48__std__lane26_strm0_data_valid  ,

            // manager 48, lane 26, stream 1      
            input   wire                                        std__mgr48__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane26_strm1_data        ,
            output  wire                                        mgr48__std__lane26_strm1_data_valid  ,

            // manager 48, lane 27, stream 0      
            input   wire                                        std__mgr48__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane27_strm0_data        ,
            output  wire                                        mgr48__std__lane27_strm0_data_valid  ,

            // manager 48, lane 27, stream 1      
            input   wire                                        std__mgr48__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane27_strm1_data        ,
            output  wire                                        mgr48__std__lane27_strm1_data_valid  ,

            // manager 48, lane 28, stream 0      
            input   wire                                        std__mgr48__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane28_strm0_data        ,
            output  wire                                        mgr48__std__lane28_strm0_data_valid  ,

            // manager 48, lane 28, stream 1      
            input   wire                                        std__mgr48__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane28_strm1_data        ,
            output  wire                                        mgr48__std__lane28_strm1_data_valid  ,

            // manager 48, lane 29, stream 0      
            input   wire                                        std__mgr48__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane29_strm0_data        ,
            output  wire                                        mgr48__std__lane29_strm0_data_valid  ,

            // manager 48, lane 29, stream 1      
            input   wire                                        std__mgr48__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane29_strm1_data        ,
            output  wire                                        mgr48__std__lane29_strm1_data_valid  ,

            // manager 48, lane 30, stream 0      
            input   wire                                        std__mgr48__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane30_strm0_data        ,
            output  wire                                        mgr48__std__lane30_strm0_data_valid  ,

            // manager 48, lane 30, stream 1      
            input   wire                                        std__mgr48__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane30_strm1_data        ,
            output  wire                                        mgr48__std__lane30_strm1_data_valid  ,

            // manager 48, lane 31, stream 0      
            input   wire                                        std__mgr48__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane31_strm0_data        ,
            output  wire                                        mgr48__std__lane31_strm0_data_valid  ,

            // manager 48, lane 31, stream 1      
            input   wire                                        std__mgr48__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr48__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr48__std__lane31_strm1_data        ,
            output  wire                                        mgr48__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 49, lane 0, stream 0      
            input   wire                                        std__mgr49__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane0_strm0_data        ,
            output  wire                                        mgr49__std__lane0_strm0_data_valid  ,

            // manager 49, lane 0, stream 1      
            input   wire                                        std__mgr49__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane0_strm1_data        ,
            output  wire                                        mgr49__std__lane0_strm1_data_valid  ,

            // manager 49, lane 1, stream 0      
            input   wire                                        std__mgr49__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane1_strm0_data        ,
            output  wire                                        mgr49__std__lane1_strm0_data_valid  ,

            // manager 49, lane 1, stream 1      
            input   wire                                        std__mgr49__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane1_strm1_data        ,
            output  wire                                        mgr49__std__lane1_strm1_data_valid  ,

            // manager 49, lane 2, stream 0      
            input   wire                                        std__mgr49__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane2_strm0_data        ,
            output  wire                                        mgr49__std__lane2_strm0_data_valid  ,

            // manager 49, lane 2, stream 1      
            input   wire                                        std__mgr49__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane2_strm1_data        ,
            output  wire                                        mgr49__std__lane2_strm1_data_valid  ,

            // manager 49, lane 3, stream 0      
            input   wire                                        std__mgr49__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane3_strm0_data        ,
            output  wire                                        mgr49__std__lane3_strm0_data_valid  ,

            // manager 49, lane 3, stream 1      
            input   wire                                        std__mgr49__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane3_strm1_data        ,
            output  wire                                        mgr49__std__lane3_strm1_data_valid  ,

            // manager 49, lane 4, stream 0      
            input   wire                                        std__mgr49__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane4_strm0_data        ,
            output  wire                                        mgr49__std__lane4_strm0_data_valid  ,

            // manager 49, lane 4, stream 1      
            input   wire                                        std__mgr49__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane4_strm1_data        ,
            output  wire                                        mgr49__std__lane4_strm1_data_valid  ,

            // manager 49, lane 5, stream 0      
            input   wire                                        std__mgr49__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane5_strm0_data        ,
            output  wire                                        mgr49__std__lane5_strm0_data_valid  ,

            // manager 49, lane 5, stream 1      
            input   wire                                        std__mgr49__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane5_strm1_data        ,
            output  wire                                        mgr49__std__lane5_strm1_data_valid  ,

            // manager 49, lane 6, stream 0      
            input   wire                                        std__mgr49__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane6_strm0_data        ,
            output  wire                                        mgr49__std__lane6_strm0_data_valid  ,

            // manager 49, lane 6, stream 1      
            input   wire                                        std__mgr49__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane6_strm1_data        ,
            output  wire                                        mgr49__std__lane6_strm1_data_valid  ,

            // manager 49, lane 7, stream 0      
            input   wire                                        std__mgr49__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane7_strm0_data        ,
            output  wire                                        mgr49__std__lane7_strm0_data_valid  ,

            // manager 49, lane 7, stream 1      
            input   wire                                        std__mgr49__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane7_strm1_data        ,
            output  wire                                        mgr49__std__lane7_strm1_data_valid  ,

            // manager 49, lane 8, stream 0      
            input   wire                                        std__mgr49__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane8_strm0_data        ,
            output  wire                                        mgr49__std__lane8_strm0_data_valid  ,

            // manager 49, lane 8, stream 1      
            input   wire                                        std__mgr49__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane8_strm1_data        ,
            output  wire                                        mgr49__std__lane8_strm1_data_valid  ,

            // manager 49, lane 9, stream 0      
            input   wire                                        std__mgr49__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane9_strm0_data        ,
            output  wire                                        mgr49__std__lane9_strm0_data_valid  ,

            // manager 49, lane 9, stream 1      
            input   wire                                        std__mgr49__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane9_strm1_data        ,
            output  wire                                        mgr49__std__lane9_strm1_data_valid  ,

            // manager 49, lane 10, stream 0      
            input   wire                                        std__mgr49__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane10_strm0_data        ,
            output  wire                                        mgr49__std__lane10_strm0_data_valid  ,

            // manager 49, lane 10, stream 1      
            input   wire                                        std__mgr49__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane10_strm1_data        ,
            output  wire                                        mgr49__std__lane10_strm1_data_valid  ,

            // manager 49, lane 11, stream 0      
            input   wire                                        std__mgr49__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane11_strm0_data        ,
            output  wire                                        mgr49__std__lane11_strm0_data_valid  ,

            // manager 49, lane 11, stream 1      
            input   wire                                        std__mgr49__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane11_strm1_data        ,
            output  wire                                        mgr49__std__lane11_strm1_data_valid  ,

            // manager 49, lane 12, stream 0      
            input   wire                                        std__mgr49__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane12_strm0_data        ,
            output  wire                                        mgr49__std__lane12_strm0_data_valid  ,

            // manager 49, lane 12, stream 1      
            input   wire                                        std__mgr49__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane12_strm1_data        ,
            output  wire                                        mgr49__std__lane12_strm1_data_valid  ,

            // manager 49, lane 13, stream 0      
            input   wire                                        std__mgr49__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane13_strm0_data        ,
            output  wire                                        mgr49__std__lane13_strm0_data_valid  ,

            // manager 49, lane 13, stream 1      
            input   wire                                        std__mgr49__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane13_strm1_data        ,
            output  wire                                        mgr49__std__lane13_strm1_data_valid  ,

            // manager 49, lane 14, stream 0      
            input   wire                                        std__mgr49__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane14_strm0_data        ,
            output  wire                                        mgr49__std__lane14_strm0_data_valid  ,

            // manager 49, lane 14, stream 1      
            input   wire                                        std__mgr49__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane14_strm1_data        ,
            output  wire                                        mgr49__std__lane14_strm1_data_valid  ,

            // manager 49, lane 15, stream 0      
            input   wire                                        std__mgr49__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane15_strm0_data        ,
            output  wire                                        mgr49__std__lane15_strm0_data_valid  ,

            // manager 49, lane 15, stream 1      
            input   wire                                        std__mgr49__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane15_strm1_data        ,
            output  wire                                        mgr49__std__lane15_strm1_data_valid  ,

            // manager 49, lane 16, stream 0      
            input   wire                                        std__mgr49__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane16_strm0_data        ,
            output  wire                                        mgr49__std__lane16_strm0_data_valid  ,

            // manager 49, lane 16, stream 1      
            input   wire                                        std__mgr49__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane16_strm1_data        ,
            output  wire                                        mgr49__std__lane16_strm1_data_valid  ,

            // manager 49, lane 17, stream 0      
            input   wire                                        std__mgr49__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane17_strm0_data        ,
            output  wire                                        mgr49__std__lane17_strm0_data_valid  ,

            // manager 49, lane 17, stream 1      
            input   wire                                        std__mgr49__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane17_strm1_data        ,
            output  wire                                        mgr49__std__lane17_strm1_data_valid  ,

            // manager 49, lane 18, stream 0      
            input   wire                                        std__mgr49__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane18_strm0_data        ,
            output  wire                                        mgr49__std__lane18_strm0_data_valid  ,

            // manager 49, lane 18, stream 1      
            input   wire                                        std__mgr49__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane18_strm1_data        ,
            output  wire                                        mgr49__std__lane18_strm1_data_valid  ,

            // manager 49, lane 19, stream 0      
            input   wire                                        std__mgr49__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane19_strm0_data        ,
            output  wire                                        mgr49__std__lane19_strm0_data_valid  ,

            // manager 49, lane 19, stream 1      
            input   wire                                        std__mgr49__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane19_strm1_data        ,
            output  wire                                        mgr49__std__lane19_strm1_data_valid  ,

            // manager 49, lane 20, stream 0      
            input   wire                                        std__mgr49__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane20_strm0_data        ,
            output  wire                                        mgr49__std__lane20_strm0_data_valid  ,

            // manager 49, lane 20, stream 1      
            input   wire                                        std__mgr49__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane20_strm1_data        ,
            output  wire                                        mgr49__std__lane20_strm1_data_valid  ,

            // manager 49, lane 21, stream 0      
            input   wire                                        std__mgr49__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane21_strm0_data        ,
            output  wire                                        mgr49__std__lane21_strm0_data_valid  ,

            // manager 49, lane 21, stream 1      
            input   wire                                        std__mgr49__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane21_strm1_data        ,
            output  wire                                        mgr49__std__lane21_strm1_data_valid  ,

            // manager 49, lane 22, stream 0      
            input   wire                                        std__mgr49__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane22_strm0_data        ,
            output  wire                                        mgr49__std__lane22_strm0_data_valid  ,

            // manager 49, lane 22, stream 1      
            input   wire                                        std__mgr49__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane22_strm1_data        ,
            output  wire                                        mgr49__std__lane22_strm1_data_valid  ,

            // manager 49, lane 23, stream 0      
            input   wire                                        std__mgr49__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane23_strm0_data        ,
            output  wire                                        mgr49__std__lane23_strm0_data_valid  ,

            // manager 49, lane 23, stream 1      
            input   wire                                        std__mgr49__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane23_strm1_data        ,
            output  wire                                        mgr49__std__lane23_strm1_data_valid  ,

            // manager 49, lane 24, stream 0      
            input   wire                                        std__mgr49__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane24_strm0_data        ,
            output  wire                                        mgr49__std__lane24_strm0_data_valid  ,

            // manager 49, lane 24, stream 1      
            input   wire                                        std__mgr49__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane24_strm1_data        ,
            output  wire                                        mgr49__std__lane24_strm1_data_valid  ,

            // manager 49, lane 25, stream 0      
            input   wire                                        std__mgr49__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane25_strm0_data        ,
            output  wire                                        mgr49__std__lane25_strm0_data_valid  ,

            // manager 49, lane 25, stream 1      
            input   wire                                        std__mgr49__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane25_strm1_data        ,
            output  wire                                        mgr49__std__lane25_strm1_data_valid  ,

            // manager 49, lane 26, stream 0      
            input   wire                                        std__mgr49__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane26_strm0_data        ,
            output  wire                                        mgr49__std__lane26_strm0_data_valid  ,

            // manager 49, lane 26, stream 1      
            input   wire                                        std__mgr49__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane26_strm1_data        ,
            output  wire                                        mgr49__std__lane26_strm1_data_valid  ,

            // manager 49, lane 27, stream 0      
            input   wire                                        std__mgr49__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane27_strm0_data        ,
            output  wire                                        mgr49__std__lane27_strm0_data_valid  ,

            // manager 49, lane 27, stream 1      
            input   wire                                        std__mgr49__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane27_strm1_data        ,
            output  wire                                        mgr49__std__lane27_strm1_data_valid  ,

            // manager 49, lane 28, stream 0      
            input   wire                                        std__mgr49__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane28_strm0_data        ,
            output  wire                                        mgr49__std__lane28_strm0_data_valid  ,

            // manager 49, lane 28, stream 1      
            input   wire                                        std__mgr49__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane28_strm1_data        ,
            output  wire                                        mgr49__std__lane28_strm1_data_valid  ,

            // manager 49, lane 29, stream 0      
            input   wire                                        std__mgr49__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane29_strm0_data        ,
            output  wire                                        mgr49__std__lane29_strm0_data_valid  ,

            // manager 49, lane 29, stream 1      
            input   wire                                        std__mgr49__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane29_strm1_data        ,
            output  wire                                        mgr49__std__lane29_strm1_data_valid  ,

            // manager 49, lane 30, stream 0      
            input   wire                                        std__mgr49__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane30_strm0_data        ,
            output  wire                                        mgr49__std__lane30_strm0_data_valid  ,

            // manager 49, lane 30, stream 1      
            input   wire                                        std__mgr49__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane30_strm1_data        ,
            output  wire                                        mgr49__std__lane30_strm1_data_valid  ,

            // manager 49, lane 31, stream 0      
            input   wire                                        std__mgr49__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane31_strm0_data        ,
            output  wire                                        mgr49__std__lane31_strm0_data_valid  ,

            // manager 49, lane 31, stream 1      
            input   wire                                        std__mgr49__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr49__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr49__std__lane31_strm1_data        ,
            output  wire                                        mgr49__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 50, lane 0, stream 0      
            input   wire                                        std__mgr50__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane0_strm0_data        ,
            output  wire                                        mgr50__std__lane0_strm0_data_valid  ,

            // manager 50, lane 0, stream 1      
            input   wire                                        std__mgr50__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane0_strm1_data        ,
            output  wire                                        mgr50__std__lane0_strm1_data_valid  ,

            // manager 50, lane 1, stream 0      
            input   wire                                        std__mgr50__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane1_strm0_data        ,
            output  wire                                        mgr50__std__lane1_strm0_data_valid  ,

            // manager 50, lane 1, stream 1      
            input   wire                                        std__mgr50__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane1_strm1_data        ,
            output  wire                                        mgr50__std__lane1_strm1_data_valid  ,

            // manager 50, lane 2, stream 0      
            input   wire                                        std__mgr50__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane2_strm0_data        ,
            output  wire                                        mgr50__std__lane2_strm0_data_valid  ,

            // manager 50, lane 2, stream 1      
            input   wire                                        std__mgr50__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane2_strm1_data        ,
            output  wire                                        mgr50__std__lane2_strm1_data_valid  ,

            // manager 50, lane 3, stream 0      
            input   wire                                        std__mgr50__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane3_strm0_data        ,
            output  wire                                        mgr50__std__lane3_strm0_data_valid  ,

            // manager 50, lane 3, stream 1      
            input   wire                                        std__mgr50__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane3_strm1_data        ,
            output  wire                                        mgr50__std__lane3_strm1_data_valid  ,

            // manager 50, lane 4, stream 0      
            input   wire                                        std__mgr50__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane4_strm0_data        ,
            output  wire                                        mgr50__std__lane4_strm0_data_valid  ,

            // manager 50, lane 4, stream 1      
            input   wire                                        std__mgr50__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane4_strm1_data        ,
            output  wire                                        mgr50__std__lane4_strm1_data_valid  ,

            // manager 50, lane 5, stream 0      
            input   wire                                        std__mgr50__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane5_strm0_data        ,
            output  wire                                        mgr50__std__lane5_strm0_data_valid  ,

            // manager 50, lane 5, stream 1      
            input   wire                                        std__mgr50__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane5_strm1_data        ,
            output  wire                                        mgr50__std__lane5_strm1_data_valid  ,

            // manager 50, lane 6, stream 0      
            input   wire                                        std__mgr50__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane6_strm0_data        ,
            output  wire                                        mgr50__std__lane6_strm0_data_valid  ,

            // manager 50, lane 6, stream 1      
            input   wire                                        std__mgr50__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane6_strm1_data        ,
            output  wire                                        mgr50__std__lane6_strm1_data_valid  ,

            // manager 50, lane 7, stream 0      
            input   wire                                        std__mgr50__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane7_strm0_data        ,
            output  wire                                        mgr50__std__lane7_strm0_data_valid  ,

            // manager 50, lane 7, stream 1      
            input   wire                                        std__mgr50__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane7_strm1_data        ,
            output  wire                                        mgr50__std__lane7_strm1_data_valid  ,

            // manager 50, lane 8, stream 0      
            input   wire                                        std__mgr50__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane8_strm0_data        ,
            output  wire                                        mgr50__std__lane8_strm0_data_valid  ,

            // manager 50, lane 8, stream 1      
            input   wire                                        std__mgr50__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane8_strm1_data        ,
            output  wire                                        mgr50__std__lane8_strm1_data_valid  ,

            // manager 50, lane 9, stream 0      
            input   wire                                        std__mgr50__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane9_strm0_data        ,
            output  wire                                        mgr50__std__lane9_strm0_data_valid  ,

            // manager 50, lane 9, stream 1      
            input   wire                                        std__mgr50__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane9_strm1_data        ,
            output  wire                                        mgr50__std__lane9_strm1_data_valid  ,

            // manager 50, lane 10, stream 0      
            input   wire                                        std__mgr50__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane10_strm0_data        ,
            output  wire                                        mgr50__std__lane10_strm0_data_valid  ,

            // manager 50, lane 10, stream 1      
            input   wire                                        std__mgr50__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane10_strm1_data        ,
            output  wire                                        mgr50__std__lane10_strm1_data_valid  ,

            // manager 50, lane 11, stream 0      
            input   wire                                        std__mgr50__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane11_strm0_data        ,
            output  wire                                        mgr50__std__lane11_strm0_data_valid  ,

            // manager 50, lane 11, stream 1      
            input   wire                                        std__mgr50__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane11_strm1_data        ,
            output  wire                                        mgr50__std__lane11_strm1_data_valid  ,

            // manager 50, lane 12, stream 0      
            input   wire                                        std__mgr50__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane12_strm0_data        ,
            output  wire                                        mgr50__std__lane12_strm0_data_valid  ,

            // manager 50, lane 12, stream 1      
            input   wire                                        std__mgr50__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane12_strm1_data        ,
            output  wire                                        mgr50__std__lane12_strm1_data_valid  ,

            // manager 50, lane 13, stream 0      
            input   wire                                        std__mgr50__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane13_strm0_data        ,
            output  wire                                        mgr50__std__lane13_strm0_data_valid  ,

            // manager 50, lane 13, stream 1      
            input   wire                                        std__mgr50__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane13_strm1_data        ,
            output  wire                                        mgr50__std__lane13_strm1_data_valid  ,

            // manager 50, lane 14, stream 0      
            input   wire                                        std__mgr50__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane14_strm0_data        ,
            output  wire                                        mgr50__std__lane14_strm0_data_valid  ,

            // manager 50, lane 14, stream 1      
            input   wire                                        std__mgr50__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane14_strm1_data        ,
            output  wire                                        mgr50__std__lane14_strm1_data_valid  ,

            // manager 50, lane 15, stream 0      
            input   wire                                        std__mgr50__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane15_strm0_data        ,
            output  wire                                        mgr50__std__lane15_strm0_data_valid  ,

            // manager 50, lane 15, stream 1      
            input   wire                                        std__mgr50__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane15_strm1_data        ,
            output  wire                                        mgr50__std__lane15_strm1_data_valid  ,

            // manager 50, lane 16, stream 0      
            input   wire                                        std__mgr50__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane16_strm0_data        ,
            output  wire                                        mgr50__std__lane16_strm0_data_valid  ,

            // manager 50, lane 16, stream 1      
            input   wire                                        std__mgr50__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane16_strm1_data        ,
            output  wire                                        mgr50__std__lane16_strm1_data_valid  ,

            // manager 50, lane 17, stream 0      
            input   wire                                        std__mgr50__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane17_strm0_data        ,
            output  wire                                        mgr50__std__lane17_strm0_data_valid  ,

            // manager 50, lane 17, stream 1      
            input   wire                                        std__mgr50__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane17_strm1_data        ,
            output  wire                                        mgr50__std__lane17_strm1_data_valid  ,

            // manager 50, lane 18, stream 0      
            input   wire                                        std__mgr50__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane18_strm0_data        ,
            output  wire                                        mgr50__std__lane18_strm0_data_valid  ,

            // manager 50, lane 18, stream 1      
            input   wire                                        std__mgr50__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane18_strm1_data        ,
            output  wire                                        mgr50__std__lane18_strm1_data_valid  ,

            // manager 50, lane 19, stream 0      
            input   wire                                        std__mgr50__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane19_strm0_data        ,
            output  wire                                        mgr50__std__lane19_strm0_data_valid  ,

            // manager 50, lane 19, stream 1      
            input   wire                                        std__mgr50__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane19_strm1_data        ,
            output  wire                                        mgr50__std__lane19_strm1_data_valid  ,

            // manager 50, lane 20, stream 0      
            input   wire                                        std__mgr50__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane20_strm0_data        ,
            output  wire                                        mgr50__std__lane20_strm0_data_valid  ,

            // manager 50, lane 20, stream 1      
            input   wire                                        std__mgr50__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane20_strm1_data        ,
            output  wire                                        mgr50__std__lane20_strm1_data_valid  ,

            // manager 50, lane 21, stream 0      
            input   wire                                        std__mgr50__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane21_strm0_data        ,
            output  wire                                        mgr50__std__lane21_strm0_data_valid  ,

            // manager 50, lane 21, stream 1      
            input   wire                                        std__mgr50__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane21_strm1_data        ,
            output  wire                                        mgr50__std__lane21_strm1_data_valid  ,

            // manager 50, lane 22, stream 0      
            input   wire                                        std__mgr50__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane22_strm0_data        ,
            output  wire                                        mgr50__std__lane22_strm0_data_valid  ,

            // manager 50, lane 22, stream 1      
            input   wire                                        std__mgr50__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane22_strm1_data        ,
            output  wire                                        mgr50__std__lane22_strm1_data_valid  ,

            // manager 50, lane 23, stream 0      
            input   wire                                        std__mgr50__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane23_strm0_data        ,
            output  wire                                        mgr50__std__lane23_strm0_data_valid  ,

            // manager 50, lane 23, stream 1      
            input   wire                                        std__mgr50__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane23_strm1_data        ,
            output  wire                                        mgr50__std__lane23_strm1_data_valid  ,

            // manager 50, lane 24, stream 0      
            input   wire                                        std__mgr50__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane24_strm0_data        ,
            output  wire                                        mgr50__std__lane24_strm0_data_valid  ,

            // manager 50, lane 24, stream 1      
            input   wire                                        std__mgr50__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane24_strm1_data        ,
            output  wire                                        mgr50__std__lane24_strm1_data_valid  ,

            // manager 50, lane 25, stream 0      
            input   wire                                        std__mgr50__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane25_strm0_data        ,
            output  wire                                        mgr50__std__lane25_strm0_data_valid  ,

            // manager 50, lane 25, stream 1      
            input   wire                                        std__mgr50__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane25_strm1_data        ,
            output  wire                                        mgr50__std__lane25_strm1_data_valid  ,

            // manager 50, lane 26, stream 0      
            input   wire                                        std__mgr50__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane26_strm0_data        ,
            output  wire                                        mgr50__std__lane26_strm0_data_valid  ,

            // manager 50, lane 26, stream 1      
            input   wire                                        std__mgr50__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane26_strm1_data        ,
            output  wire                                        mgr50__std__lane26_strm1_data_valid  ,

            // manager 50, lane 27, stream 0      
            input   wire                                        std__mgr50__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane27_strm0_data        ,
            output  wire                                        mgr50__std__lane27_strm0_data_valid  ,

            // manager 50, lane 27, stream 1      
            input   wire                                        std__mgr50__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane27_strm1_data        ,
            output  wire                                        mgr50__std__lane27_strm1_data_valid  ,

            // manager 50, lane 28, stream 0      
            input   wire                                        std__mgr50__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane28_strm0_data        ,
            output  wire                                        mgr50__std__lane28_strm0_data_valid  ,

            // manager 50, lane 28, stream 1      
            input   wire                                        std__mgr50__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane28_strm1_data        ,
            output  wire                                        mgr50__std__lane28_strm1_data_valid  ,

            // manager 50, lane 29, stream 0      
            input   wire                                        std__mgr50__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane29_strm0_data        ,
            output  wire                                        mgr50__std__lane29_strm0_data_valid  ,

            // manager 50, lane 29, stream 1      
            input   wire                                        std__mgr50__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane29_strm1_data        ,
            output  wire                                        mgr50__std__lane29_strm1_data_valid  ,

            // manager 50, lane 30, stream 0      
            input   wire                                        std__mgr50__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane30_strm0_data        ,
            output  wire                                        mgr50__std__lane30_strm0_data_valid  ,

            // manager 50, lane 30, stream 1      
            input   wire                                        std__mgr50__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane30_strm1_data        ,
            output  wire                                        mgr50__std__lane30_strm1_data_valid  ,

            // manager 50, lane 31, stream 0      
            input   wire                                        std__mgr50__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane31_strm0_data        ,
            output  wire                                        mgr50__std__lane31_strm0_data_valid  ,

            // manager 50, lane 31, stream 1      
            input   wire                                        std__mgr50__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr50__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr50__std__lane31_strm1_data        ,
            output  wire                                        mgr50__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 51, lane 0, stream 0      
            input   wire                                        std__mgr51__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane0_strm0_data        ,
            output  wire                                        mgr51__std__lane0_strm0_data_valid  ,

            // manager 51, lane 0, stream 1      
            input   wire                                        std__mgr51__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane0_strm1_data        ,
            output  wire                                        mgr51__std__lane0_strm1_data_valid  ,

            // manager 51, lane 1, stream 0      
            input   wire                                        std__mgr51__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane1_strm0_data        ,
            output  wire                                        mgr51__std__lane1_strm0_data_valid  ,

            // manager 51, lane 1, stream 1      
            input   wire                                        std__mgr51__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane1_strm1_data        ,
            output  wire                                        mgr51__std__lane1_strm1_data_valid  ,

            // manager 51, lane 2, stream 0      
            input   wire                                        std__mgr51__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane2_strm0_data        ,
            output  wire                                        mgr51__std__lane2_strm0_data_valid  ,

            // manager 51, lane 2, stream 1      
            input   wire                                        std__mgr51__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane2_strm1_data        ,
            output  wire                                        mgr51__std__lane2_strm1_data_valid  ,

            // manager 51, lane 3, stream 0      
            input   wire                                        std__mgr51__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane3_strm0_data        ,
            output  wire                                        mgr51__std__lane3_strm0_data_valid  ,

            // manager 51, lane 3, stream 1      
            input   wire                                        std__mgr51__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane3_strm1_data        ,
            output  wire                                        mgr51__std__lane3_strm1_data_valid  ,

            // manager 51, lane 4, stream 0      
            input   wire                                        std__mgr51__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane4_strm0_data        ,
            output  wire                                        mgr51__std__lane4_strm0_data_valid  ,

            // manager 51, lane 4, stream 1      
            input   wire                                        std__mgr51__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane4_strm1_data        ,
            output  wire                                        mgr51__std__lane4_strm1_data_valid  ,

            // manager 51, lane 5, stream 0      
            input   wire                                        std__mgr51__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane5_strm0_data        ,
            output  wire                                        mgr51__std__lane5_strm0_data_valid  ,

            // manager 51, lane 5, stream 1      
            input   wire                                        std__mgr51__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane5_strm1_data        ,
            output  wire                                        mgr51__std__lane5_strm1_data_valid  ,

            // manager 51, lane 6, stream 0      
            input   wire                                        std__mgr51__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane6_strm0_data        ,
            output  wire                                        mgr51__std__lane6_strm0_data_valid  ,

            // manager 51, lane 6, stream 1      
            input   wire                                        std__mgr51__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane6_strm1_data        ,
            output  wire                                        mgr51__std__lane6_strm1_data_valid  ,

            // manager 51, lane 7, stream 0      
            input   wire                                        std__mgr51__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane7_strm0_data        ,
            output  wire                                        mgr51__std__lane7_strm0_data_valid  ,

            // manager 51, lane 7, stream 1      
            input   wire                                        std__mgr51__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane7_strm1_data        ,
            output  wire                                        mgr51__std__lane7_strm1_data_valid  ,

            // manager 51, lane 8, stream 0      
            input   wire                                        std__mgr51__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane8_strm0_data        ,
            output  wire                                        mgr51__std__lane8_strm0_data_valid  ,

            // manager 51, lane 8, stream 1      
            input   wire                                        std__mgr51__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane8_strm1_data        ,
            output  wire                                        mgr51__std__lane8_strm1_data_valid  ,

            // manager 51, lane 9, stream 0      
            input   wire                                        std__mgr51__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane9_strm0_data        ,
            output  wire                                        mgr51__std__lane9_strm0_data_valid  ,

            // manager 51, lane 9, stream 1      
            input   wire                                        std__mgr51__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane9_strm1_data        ,
            output  wire                                        mgr51__std__lane9_strm1_data_valid  ,

            // manager 51, lane 10, stream 0      
            input   wire                                        std__mgr51__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane10_strm0_data        ,
            output  wire                                        mgr51__std__lane10_strm0_data_valid  ,

            // manager 51, lane 10, stream 1      
            input   wire                                        std__mgr51__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane10_strm1_data        ,
            output  wire                                        mgr51__std__lane10_strm1_data_valid  ,

            // manager 51, lane 11, stream 0      
            input   wire                                        std__mgr51__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane11_strm0_data        ,
            output  wire                                        mgr51__std__lane11_strm0_data_valid  ,

            // manager 51, lane 11, stream 1      
            input   wire                                        std__mgr51__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane11_strm1_data        ,
            output  wire                                        mgr51__std__lane11_strm1_data_valid  ,

            // manager 51, lane 12, stream 0      
            input   wire                                        std__mgr51__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane12_strm0_data        ,
            output  wire                                        mgr51__std__lane12_strm0_data_valid  ,

            // manager 51, lane 12, stream 1      
            input   wire                                        std__mgr51__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane12_strm1_data        ,
            output  wire                                        mgr51__std__lane12_strm1_data_valid  ,

            // manager 51, lane 13, stream 0      
            input   wire                                        std__mgr51__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane13_strm0_data        ,
            output  wire                                        mgr51__std__lane13_strm0_data_valid  ,

            // manager 51, lane 13, stream 1      
            input   wire                                        std__mgr51__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane13_strm1_data        ,
            output  wire                                        mgr51__std__lane13_strm1_data_valid  ,

            // manager 51, lane 14, stream 0      
            input   wire                                        std__mgr51__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane14_strm0_data        ,
            output  wire                                        mgr51__std__lane14_strm0_data_valid  ,

            // manager 51, lane 14, stream 1      
            input   wire                                        std__mgr51__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane14_strm1_data        ,
            output  wire                                        mgr51__std__lane14_strm1_data_valid  ,

            // manager 51, lane 15, stream 0      
            input   wire                                        std__mgr51__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane15_strm0_data        ,
            output  wire                                        mgr51__std__lane15_strm0_data_valid  ,

            // manager 51, lane 15, stream 1      
            input   wire                                        std__mgr51__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane15_strm1_data        ,
            output  wire                                        mgr51__std__lane15_strm1_data_valid  ,

            // manager 51, lane 16, stream 0      
            input   wire                                        std__mgr51__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane16_strm0_data        ,
            output  wire                                        mgr51__std__lane16_strm0_data_valid  ,

            // manager 51, lane 16, stream 1      
            input   wire                                        std__mgr51__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane16_strm1_data        ,
            output  wire                                        mgr51__std__lane16_strm1_data_valid  ,

            // manager 51, lane 17, stream 0      
            input   wire                                        std__mgr51__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane17_strm0_data        ,
            output  wire                                        mgr51__std__lane17_strm0_data_valid  ,

            // manager 51, lane 17, stream 1      
            input   wire                                        std__mgr51__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane17_strm1_data        ,
            output  wire                                        mgr51__std__lane17_strm1_data_valid  ,

            // manager 51, lane 18, stream 0      
            input   wire                                        std__mgr51__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane18_strm0_data        ,
            output  wire                                        mgr51__std__lane18_strm0_data_valid  ,

            // manager 51, lane 18, stream 1      
            input   wire                                        std__mgr51__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane18_strm1_data        ,
            output  wire                                        mgr51__std__lane18_strm1_data_valid  ,

            // manager 51, lane 19, stream 0      
            input   wire                                        std__mgr51__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane19_strm0_data        ,
            output  wire                                        mgr51__std__lane19_strm0_data_valid  ,

            // manager 51, lane 19, stream 1      
            input   wire                                        std__mgr51__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane19_strm1_data        ,
            output  wire                                        mgr51__std__lane19_strm1_data_valid  ,

            // manager 51, lane 20, stream 0      
            input   wire                                        std__mgr51__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane20_strm0_data        ,
            output  wire                                        mgr51__std__lane20_strm0_data_valid  ,

            // manager 51, lane 20, stream 1      
            input   wire                                        std__mgr51__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane20_strm1_data        ,
            output  wire                                        mgr51__std__lane20_strm1_data_valid  ,

            // manager 51, lane 21, stream 0      
            input   wire                                        std__mgr51__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane21_strm0_data        ,
            output  wire                                        mgr51__std__lane21_strm0_data_valid  ,

            // manager 51, lane 21, stream 1      
            input   wire                                        std__mgr51__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane21_strm1_data        ,
            output  wire                                        mgr51__std__lane21_strm1_data_valid  ,

            // manager 51, lane 22, stream 0      
            input   wire                                        std__mgr51__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane22_strm0_data        ,
            output  wire                                        mgr51__std__lane22_strm0_data_valid  ,

            // manager 51, lane 22, stream 1      
            input   wire                                        std__mgr51__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane22_strm1_data        ,
            output  wire                                        mgr51__std__lane22_strm1_data_valid  ,

            // manager 51, lane 23, stream 0      
            input   wire                                        std__mgr51__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane23_strm0_data        ,
            output  wire                                        mgr51__std__lane23_strm0_data_valid  ,

            // manager 51, lane 23, stream 1      
            input   wire                                        std__mgr51__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane23_strm1_data        ,
            output  wire                                        mgr51__std__lane23_strm1_data_valid  ,

            // manager 51, lane 24, stream 0      
            input   wire                                        std__mgr51__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane24_strm0_data        ,
            output  wire                                        mgr51__std__lane24_strm0_data_valid  ,

            // manager 51, lane 24, stream 1      
            input   wire                                        std__mgr51__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane24_strm1_data        ,
            output  wire                                        mgr51__std__lane24_strm1_data_valid  ,

            // manager 51, lane 25, stream 0      
            input   wire                                        std__mgr51__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane25_strm0_data        ,
            output  wire                                        mgr51__std__lane25_strm0_data_valid  ,

            // manager 51, lane 25, stream 1      
            input   wire                                        std__mgr51__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane25_strm1_data        ,
            output  wire                                        mgr51__std__lane25_strm1_data_valid  ,

            // manager 51, lane 26, stream 0      
            input   wire                                        std__mgr51__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane26_strm0_data        ,
            output  wire                                        mgr51__std__lane26_strm0_data_valid  ,

            // manager 51, lane 26, stream 1      
            input   wire                                        std__mgr51__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane26_strm1_data        ,
            output  wire                                        mgr51__std__lane26_strm1_data_valid  ,

            // manager 51, lane 27, stream 0      
            input   wire                                        std__mgr51__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane27_strm0_data        ,
            output  wire                                        mgr51__std__lane27_strm0_data_valid  ,

            // manager 51, lane 27, stream 1      
            input   wire                                        std__mgr51__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane27_strm1_data        ,
            output  wire                                        mgr51__std__lane27_strm1_data_valid  ,

            // manager 51, lane 28, stream 0      
            input   wire                                        std__mgr51__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane28_strm0_data        ,
            output  wire                                        mgr51__std__lane28_strm0_data_valid  ,

            // manager 51, lane 28, stream 1      
            input   wire                                        std__mgr51__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane28_strm1_data        ,
            output  wire                                        mgr51__std__lane28_strm1_data_valid  ,

            // manager 51, lane 29, stream 0      
            input   wire                                        std__mgr51__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane29_strm0_data        ,
            output  wire                                        mgr51__std__lane29_strm0_data_valid  ,

            // manager 51, lane 29, stream 1      
            input   wire                                        std__mgr51__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane29_strm1_data        ,
            output  wire                                        mgr51__std__lane29_strm1_data_valid  ,

            // manager 51, lane 30, stream 0      
            input   wire                                        std__mgr51__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane30_strm0_data        ,
            output  wire                                        mgr51__std__lane30_strm0_data_valid  ,

            // manager 51, lane 30, stream 1      
            input   wire                                        std__mgr51__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane30_strm1_data        ,
            output  wire                                        mgr51__std__lane30_strm1_data_valid  ,

            // manager 51, lane 31, stream 0      
            input   wire                                        std__mgr51__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane31_strm0_data        ,
            output  wire                                        mgr51__std__lane31_strm0_data_valid  ,

            // manager 51, lane 31, stream 1      
            input   wire                                        std__mgr51__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr51__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr51__std__lane31_strm1_data        ,
            output  wire                                        mgr51__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 52, lane 0, stream 0      
            input   wire                                        std__mgr52__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane0_strm0_data        ,
            output  wire                                        mgr52__std__lane0_strm0_data_valid  ,

            // manager 52, lane 0, stream 1      
            input   wire                                        std__mgr52__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane0_strm1_data        ,
            output  wire                                        mgr52__std__lane0_strm1_data_valid  ,

            // manager 52, lane 1, stream 0      
            input   wire                                        std__mgr52__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane1_strm0_data        ,
            output  wire                                        mgr52__std__lane1_strm0_data_valid  ,

            // manager 52, lane 1, stream 1      
            input   wire                                        std__mgr52__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane1_strm1_data        ,
            output  wire                                        mgr52__std__lane1_strm1_data_valid  ,

            // manager 52, lane 2, stream 0      
            input   wire                                        std__mgr52__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane2_strm0_data        ,
            output  wire                                        mgr52__std__lane2_strm0_data_valid  ,

            // manager 52, lane 2, stream 1      
            input   wire                                        std__mgr52__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane2_strm1_data        ,
            output  wire                                        mgr52__std__lane2_strm1_data_valid  ,

            // manager 52, lane 3, stream 0      
            input   wire                                        std__mgr52__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane3_strm0_data        ,
            output  wire                                        mgr52__std__lane3_strm0_data_valid  ,

            // manager 52, lane 3, stream 1      
            input   wire                                        std__mgr52__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane3_strm1_data        ,
            output  wire                                        mgr52__std__lane3_strm1_data_valid  ,

            // manager 52, lane 4, stream 0      
            input   wire                                        std__mgr52__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane4_strm0_data        ,
            output  wire                                        mgr52__std__lane4_strm0_data_valid  ,

            // manager 52, lane 4, stream 1      
            input   wire                                        std__mgr52__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane4_strm1_data        ,
            output  wire                                        mgr52__std__lane4_strm1_data_valid  ,

            // manager 52, lane 5, stream 0      
            input   wire                                        std__mgr52__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane5_strm0_data        ,
            output  wire                                        mgr52__std__lane5_strm0_data_valid  ,

            // manager 52, lane 5, stream 1      
            input   wire                                        std__mgr52__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane5_strm1_data        ,
            output  wire                                        mgr52__std__lane5_strm1_data_valid  ,

            // manager 52, lane 6, stream 0      
            input   wire                                        std__mgr52__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane6_strm0_data        ,
            output  wire                                        mgr52__std__lane6_strm0_data_valid  ,

            // manager 52, lane 6, stream 1      
            input   wire                                        std__mgr52__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane6_strm1_data        ,
            output  wire                                        mgr52__std__lane6_strm1_data_valid  ,

            // manager 52, lane 7, stream 0      
            input   wire                                        std__mgr52__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane7_strm0_data        ,
            output  wire                                        mgr52__std__lane7_strm0_data_valid  ,

            // manager 52, lane 7, stream 1      
            input   wire                                        std__mgr52__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane7_strm1_data        ,
            output  wire                                        mgr52__std__lane7_strm1_data_valid  ,

            // manager 52, lane 8, stream 0      
            input   wire                                        std__mgr52__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane8_strm0_data        ,
            output  wire                                        mgr52__std__lane8_strm0_data_valid  ,

            // manager 52, lane 8, stream 1      
            input   wire                                        std__mgr52__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane8_strm1_data        ,
            output  wire                                        mgr52__std__lane8_strm1_data_valid  ,

            // manager 52, lane 9, stream 0      
            input   wire                                        std__mgr52__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane9_strm0_data        ,
            output  wire                                        mgr52__std__lane9_strm0_data_valid  ,

            // manager 52, lane 9, stream 1      
            input   wire                                        std__mgr52__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane9_strm1_data        ,
            output  wire                                        mgr52__std__lane9_strm1_data_valid  ,

            // manager 52, lane 10, stream 0      
            input   wire                                        std__mgr52__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane10_strm0_data        ,
            output  wire                                        mgr52__std__lane10_strm0_data_valid  ,

            // manager 52, lane 10, stream 1      
            input   wire                                        std__mgr52__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane10_strm1_data        ,
            output  wire                                        mgr52__std__lane10_strm1_data_valid  ,

            // manager 52, lane 11, stream 0      
            input   wire                                        std__mgr52__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane11_strm0_data        ,
            output  wire                                        mgr52__std__lane11_strm0_data_valid  ,

            // manager 52, lane 11, stream 1      
            input   wire                                        std__mgr52__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane11_strm1_data        ,
            output  wire                                        mgr52__std__lane11_strm1_data_valid  ,

            // manager 52, lane 12, stream 0      
            input   wire                                        std__mgr52__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane12_strm0_data        ,
            output  wire                                        mgr52__std__lane12_strm0_data_valid  ,

            // manager 52, lane 12, stream 1      
            input   wire                                        std__mgr52__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane12_strm1_data        ,
            output  wire                                        mgr52__std__lane12_strm1_data_valid  ,

            // manager 52, lane 13, stream 0      
            input   wire                                        std__mgr52__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane13_strm0_data        ,
            output  wire                                        mgr52__std__lane13_strm0_data_valid  ,

            // manager 52, lane 13, stream 1      
            input   wire                                        std__mgr52__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane13_strm1_data        ,
            output  wire                                        mgr52__std__lane13_strm1_data_valid  ,

            // manager 52, lane 14, stream 0      
            input   wire                                        std__mgr52__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane14_strm0_data        ,
            output  wire                                        mgr52__std__lane14_strm0_data_valid  ,

            // manager 52, lane 14, stream 1      
            input   wire                                        std__mgr52__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane14_strm1_data        ,
            output  wire                                        mgr52__std__lane14_strm1_data_valid  ,

            // manager 52, lane 15, stream 0      
            input   wire                                        std__mgr52__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane15_strm0_data        ,
            output  wire                                        mgr52__std__lane15_strm0_data_valid  ,

            // manager 52, lane 15, stream 1      
            input   wire                                        std__mgr52__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane15_strm1_data        ,
            output  wire                                        mgr52__std__lane15_strm1_data_valid  ,

            // manager 52, lane 16, stream 0      
            input   wire                                        std__mgr52__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane16_strm0_data        ,
            output  wire                                        mgr52__std__lane16_strm0_data_valid  ,

            // manager 52, lane 16, stream 1      
            input   wire                                        std__mgr52__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane16_strm1_data        ,
            output  wire                                        mgr52__std__lane16_strm1_data_valid  ,

            // manager 52, lane 17, stream 0      
            input   wire                                        std__mgr52__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane17_strm0_data        ,
            output  wire                                        mgr52__std__lane17_strm0_data_valid  ,

            // manager 52, lane 17, stream 1      
            input   wire                                        std__mgr52__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane17_strm1_data        ,
            output  wire                                        mgr52__std__lane17_strm1_data_valid  ,

            // manager 52, lane 18, stream 0      
            input   wire                                        std__mgr52__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane18_strm0_data        ,
            output  wire                                        mgr52__std__lane18_strm0_data_valid  ,

            // manager 52, lane 18, stream 1      
            input   wire                                        std__mgr52__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane18_strm1_data        ,
            output  wire                                        mgr52__std__lane18_strm1_data_valid  ,

            // manager 52, lane 19, stream 0      
            input   wire                                        std__mgr52__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane19_strm0_data        ,
            output  wire                                        mgr52__std__lane19_strm0_data_valid  ,

            // manager 52, lane 19, stream 1      
            input   wire                                        std__mgr52__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane19_strm1_data        ,
            output  wire                                        mgr52__std__lane19_strm1_data_valid  ,

            // manager 52, lane 20, stream 0      
            input   wire                                        std__mgr52__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane20_strm0_data        ,
            output  wire                                        mgr52__std__lane20_strm0_data_valid  ,

            // manager 52, lane 20, stream 1      
            input   wire                                        std__mgr52__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane20_strm1_data        ,
            output  wire                                        mgr52__std__lane20_strm1_data_valid  ,

            // manager 52, lane 21, stream 0      
            input   wire                                        std__mgr52__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane21_strm0_data        ,
            output  wire                                        mgr52__std__lane21_strm0_data_valid  ,

            // manager 52, lane 21, stream 1      
            input   wire                                        std__mgr52__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane21_strm1_data        ,
            output  wire                                        mgr52__std__lane21_strm1_data_valid  ,

            // manager 52, lane 22, stream 0      
            input   wire                                        std__mgr52__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane22_strm0_data        ,
            output  wire                                        mgr52__std__lane22_strm0_data_valid  ,

            // manager 52, lane 22, stream 1      
            input   wire                                        std__mgr52__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane22_strm1_data        ,
            output  wire                                        mgr52__std__lane22_strm1_data_valid  ,

            // manager 52, lane 23, stream 0      
            input   wire                                        std__mgr52__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane23_strm0_data        ,
            output  wire                                        mgr52__std__lane23_strm0_data_valid  ,

            // manager 52, lane 23, stream 1      
            input   wire                                        std__mgr52__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane23_strm1_data        ,
            output  wire                                        mgr52__std__lane23_strm1_data_valid  ,

            // manager 52, lane 24, stream 0      
            input   wire                                        std__mgr52__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane24_strm0_data        ,
            output  wire                                        mgr52__std__lane24_strm0_data_valid  ,

            // manager 52, lane 24, stream 1      
            input   wire                                        std__mgr52__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane24_strm1_data        ,
            output  wire                                        mgr52__std__lane24_strm1_data_valid  ,

            // manager 52, lane 25, stream 0      
            input   wire                                        std__mgr52__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane25_strm0_data        ,
            output  wire                                        mgr52__std__lane25_strm0_data_valid  ,

            // manager 52, lane 25, stream 1      
            input   wire                                        std__mgr52__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane25_strm1_data        ,
            output  wire                                        mgr52__std__lane25_strm1_data_valid  ,

            // manager 52, lane 26, stream 0      
            input   wire                                        std__mgr52__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane26_strm0_data        ,
            output  wire                                        mgr52__std__lane26_strm0_data_valid  ,

            // manager 52, lane 26, stream 1      
            input   wire                                        std__mgr52__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane26_strm1_data        ,
            output  wire                                        mgr52__std__lane26_strm1_data_valid  ,

            // manager 52, lane 27, stream 0      
            input   wire                                        std__mgr52__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane27_strm0_data        ,
            output  wire                                        mgr52__std__lane27_strm0_data_valid  ,

            // manager 52, lane 27, stream 1      
            input   wire                                        std__mgr52__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane27_strm1_data        ,
            output  wire                                        mgr52__std__lane27_strm1_data_valid  ,

            // manager 52, lane 28, stream 0      
            input   wire                                        std__mgr52__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane28_strm0_data        ,
            output  wire                                        mgr52__std__lane28_strm0_data_valid  ,

            // manager 52, lane 28, stream 1      
            input   wire                                        std__mgr52__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane28_strm1_data        ,
            output  wire                                        mgr52__std__lane28_strm1_data_valid  ,

            // manager 52, lane 29, stream 0      
            input   wire                                        std__mgr52__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane29_strm0_data        ,
            output  wire                                        mgr52__std__lane29_strm0_data_valid  ,

            // manager 52, lane 29, stream 1      
            input   wire                                        std__mgr52__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane29_strm1_data        ,
            output  wire                                        mgr52__std__lane29_strm1_data_valid  ,

            // manager 52, lane 30, stream 0      
            input   wire                                        std__mgr52__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane30_strm0_data        ,
            output  wire                                        mgr52__std__lane30_strm0_data_valid  ,

            // manager 52, lane 30, stream 1      
            input   wire                                        std__mgr52__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane30_strm1_data        ,
            output  wire                                        mgr52__std__lane30_strm1_data_valid  ,

            // manager 52, lane 31, stream 0      
            input   wire                                        std__mgr52__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane31_strm0_data        ,
            output  wire                                        mgr52__std__lane31_strm0_data_valid  ,

            // manager 52, lane 31, stream 1      
            input   wire                                        std__mgr52__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr52__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr52__std__lane31_strm1_data        ,
            output  wire                                        mgr52__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 53, lane 0, stream 0      
            input   wire                                        std__mgr53__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane0_strm0_data        ,
            output  wire                                        mgr53__std__lane0_strm0_data_valid  ,

            // manager 53, lane 0, stream 1      
            input   wire                                        std__mgr53__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane0_strm1_data        ,
            output  wire                                        mgr53__std__lane0_strm1_data_valid  ,

            // manager 53, lane 1, stream 0      
            input   wire                                        std__mgr53__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane1_strm0_data        ,
            output  wire                                        mgr53__std__lane1_strm0_data_valid  ,

            // manager 53, lane 1, stream 1      
            input   wire                                        std__mgr53__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane1_strm1_data        ,
            output  wire                                        mgr53__std__lane1_strm1_data_valid  ,

            // manager 53, lane 2, stream 0      
            input   wire                                        std__mgr53__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane2_strm0_data        ,
            output  wire                                        mgr53__std__lane2_strm0_data_valid  ,

            // manager 53, lane 2, stream 1      
            input   wire                                        std__mgr53__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane2_strm1_data        ,
            output  wire                                        mgr53__std__lane2_strm1_data_valid  ,

            // manager 53, lane 3, stream 0      
            input   wire                                        std__mgr53__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane3_strm0_data        ,
            output  wire                                        mgr53__std__lane3_strm0_data_valid  ,

            // manager 53, lane 3, stream 1      
            input   wire                                        std__mgr53__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane3_strm1_data        ,
            output  wire                                        mgr53__std__lane3_strm1_data_valid  ,

            // manager 53, lane 4, stream 0      
            input   wire                                        std__mgr53__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane4_strm0_data        ,
            output  wire                                        mgr53__std__lane4_strm0_data_valid  ,

            // manager 53, lane 4, stream 1      
            input   wire                                        std__mgr53__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane4_strm1_data        ,
            output  wire                                        mgr53__std__lane4_strm1_data_valid  ,

            // manager 53, lane 5, stream 0      
            input   wire                                        std__mgr53__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane5_strm0_data        ,
            output  wire                                        mgr53__std__lane5_strm0_data_valid  ,

            // manager 53, lane 5, stream 1      
            input   wire                                        std__mgr53__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane5_strm1_data        ,
            output  wire                                        mgr53__std__lane5_strm1_data_valid  ,

            // manager 53, lane 6, stream 0      
            input   wire                                        std__mgr53__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane6_strm0_data        ,
            output  wire                                        mgr53__std__lane6_strm0_data_valid  ,

            // manager 53, lane 6, stream 1      
            input   wire                                        std__mgr53__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane6_strm1_data        ,
            output  wire                                        mgr53__std__lane6_strm1_data_valid  ,

            // manager 53, lane 7, stream 0      
            input   wire                                        std__mgr53__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane7_strm0_data        ,
            output  wire                                        mgr53__std__lane7_strm0_data_valid  ,

            // manager 53, lane 7, stream 1      
            input   wire                                        std__mgr53__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane7_strm1_data        ,
            output  wire                                        mgr53__std__lane7_strm1_data_valid  ,

            // manager 53, lane 8, stream 0      
            input   wire                                        std__mgr53__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane8_strm0_data        ,
            output  wire                                        mgr53__std__lane8_strm0_data_valid  ,

            // manager 53, lane 8, stream 1      
            input   wire                                        std__mgr53__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane8_strm1_data        ,
            output  wire                                        mgr53__std__lane8_strm1_data_valid  ,

            // manager 53, lane 9, stream 0      
            input   wire                                        std__mgr53__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane9_strm0_data        ,
            output  wire                                        mgr53__std__lane9_strm0_data_valid  ,

            // manager 53, lane 9, stream 1      
            input   wire                                        std__mgr53__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane9_strm1_data        ,
            output  wire                                        mgr53__std__lane9_strm1_data_valid  ,

            // manager 53, lane 10, stream 0      
            input   wire                                        std__mgr53__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane10_strm0_data        ,
            output  wire                                        mgr53__std__lane10_strm0_data_valid  ,

            // manager 53, lane 10, stream 1      
            input   wire                                        std__mgr53__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane10_strm1_data        ,
            output  wire                                        mgr53__std__lane10_strm1_data_valid  ,

            // manager 53, lane 11, stream 0      
            input   wire                                        std__mgr53__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane11_strm0_data        ,
            output  wire                                        mgr53__std__lane11_strm0_data_valid  ,

            // manager 53, lane 11, stream 1      
            input   wire                                        std__mgr53__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane11_strm1_data        ,
            output  wire                                        mgr53__std__lane11_strm1_data_valid  ,

            // manager 53, lane 12, stream 0      
            input   wire                                        std__mgr53__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane12_strm0_data        ,
            output  wire                                        mgr53__std__lane12_strm0_data_valid  ,

            // manager 53, lane 12, stream 1      
            input   wire                                        std__mgr53__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane12_strm1_data        ,
            output  wire                                        mgr53__std__lane12_strm1_data_valid  ,

            // manager 53, lane 13, stream 0      
            input   wire                                        std__mgr53__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane13_strm0_data        ,
            output  wire                                        mgr53__std__lane13_strm0_data_valid  ,

            // manager 53, lane 13, stream 1      
            input   wire                                        std__mgr53__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane13_strm1_data        ,
            output  wire                                        mgr53__std__lane13_strm1_data_valid  ,

            // manager 53, lane 14, stream 0      
            input   wire                                        std__mgr53__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane14_strm0_data        ,
            output  wire                                        mgr53__std__lane14_strm0_data_valid  ,

            // manager 53, lane 14, stream 1      
            input   wire                                        std__mgr53__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane14_strm1_data        ,
            output  wire                                        mgr53__std__lane14_strm1_data_valid  ,

            // manager 53, lane 15, stream 0      
            input   wire                                        std__mgr53__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane15_strm0_data        ,
            output  wire                                        mgr53__std__lane15_strm0_data_valid  ,

            // manager 53, lane 15, stream 1      
            input   wire                                        std__mgr53__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane15_strm1_data        ,
            output  wire                                        mgr53__std__lane15_strm1_data_valid  ,

            // manager 53, lane 16, stream 0      
            input   wire                                        std__mgr53__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane16_strm0_data        ,
            output  wire                                        mgr53__std__lane16_strm0_data_valid  ,

            // manager 53, lane 16, stream 1      
            input   wire                                        std__mgr53__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane16_strm1_data        ,
            output  wire                                        mgr53__std__lane16_strm1_data_valid  ,

            // manager 53, lane 17, stream 0      
            input   wire                                        std__mgr53__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane17_strm0_data        ,
            output  wire                                        mgr53__std__lane17_strm0_data_valid  ,

            // manager 53, lane 17, stream 1      
            input   wire                                        std__mgr53__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane17_strm1_data        ,
            output  wire                                        mgr53__std__lane17_strm1_data_valid  ,

            // manager 53, lane 18, stream 0      
            input   wire                                        std__mgr53__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane18_strm0_data        ,
            output  wire                                        mgr53__std__lane18_strm0_data_valid  ,

            // manager 53, lane 18, stream 1      
            input   wire                                        std__mgr53__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane18_strm1_data        ,
            output  wire                                        mgr53__std__lane18_strm1_data_valid  ,

            // manager 53, lane 19, stream 0      
            input   wire                                        std__mgr53__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane19_strm0_data        ,
            output  wire                                        mgr53__std__lane19_strm0_data_valid  ,

            // manager 53, lane 19, stream 1      
            input   wire                                        std__mgr53__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane19_strm1_data        ,
            output  wire                                        mgr53__std__lane19_strm1_data_valid  ,

            // manager 53, lane 20, stream 0      
            input   wire                                        std__mgr53__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane20_strm0_data        ,
            output  wire                                        mgr53__std__lane20_strm0_data_valid  ,

            // manager 53, lane 20, stream 1      
            input   wire                                        std__mgr53__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane20_strm1_data        ,
            output  wire                                        mgr53__std__lane20_strm1_data_valid  ,

            // manager 53, lane 21, stream 0      
            input   wire                                        std__mgr53__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane21_strm0_data        ,
            output  wire                                        mgr53__std__lane21_strm0_data_valid  ,

            // manager 53, lane 21, stream 1      
            input   wire                                        std__mgr53__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane21_strm1_data        ,
            output  wire                                        mgr53__std__lane21_strm1_data_valid  ,

            // manager 53, lane 22, stream 0      
            input   wire                                        std__mgr53__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane22_strm0_data        ,
            output  wire                                        mgr53__std__lane22_strm0_data_valid  ,

            // manager 53, lane 22, stream 1      
            input   wire                                        std__mgr53__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane22_strm1_data        ,
            output  wire                                        mgr53__std__lane22_strm1_data_valid  ,

            // manager 53, lane 23, stream 0      
            input   wire                                        std__mgr53__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane23_strm0_data        ,
            output  wire                                        mgr53__std__lane23_strm0_data_valid  ,

            // manager 53, lane 23, stream 1      
            input   wire                                        std__mgr53__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane23_strm1_data        ,
            output  wire                                        mgr53__std__lane23_strm1_data_valid  ,

            // manager 53, lane 24, stream 0      
            input   wire                                        std__mgr53__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane24_strm0_data        ,
            output  wire                                        mgr53__std__lane24_strm0_data_valid  ,

            // manager 53, lane 24, stream 1      
            input   wire                                        std__mgr53__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane24_strm1_data        ,
            output  wire                                        mgr53__std__lane24_strm1_data_valid  ,

            // manager 53, lane 25, stream 0      
            input   wire                                        std__mgr53__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane25_strm0_data        ,
            output  wire                                        mgr53__std__lane25_strm0_data_valid  ,

            // manager 53, lane 25, stream 1      
            input   wire                                        std__mgr53__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane25_strm1_data        ,
            output  wire                                        mgr53__std__lane25_strm1_data_valid  ,

            // manager 53, lane 26, stream 0      
            input   wire                                        std__mgr53__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane26_strm0_data        ,
            output  wire                                        mgr53__std__lane26_strm0_data_valid  ,

            // manager 53, lane 26, stream 1      
            input   wire                                        std__mgr53__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane26_strm1_data        ,
            output  wire                                        mgr53__std__lane26_strm1_data_valid  ,

            // manager 53, lane 27, stream 0      
            input   wire                                        std__mgr53__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane27_strm0_data        ,
            output  wire                                        mgr53__std__lane27_strm0_data_valid  ,

            // manager 53, lane 27, stream 1      
            input   wire                                        std__mgr53__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane27_strm1_data        ,
            output  wire                                        mgr53__std__lane27_strm1_data_valid  ,

            // manager 53, lane 28, stream 0      
            input   wire                                        std__mgr53__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane28_strm0_data        ,
            output  wire                                        mgr53__std__lane28_strm0_data_valid  ,

            // manager 53, lane 28, stream 1      
            input   wire                                        std__mgr53__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane28_strm1_data        ,
            output  wire                                        mgr53__std__lane28_strm1_data_valid  ,

            // manager 53, lane 29, stream 0      
            input   wire                                        std__mgr53__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane29_strm0_data        ,
            output  wire                                        mgr53__std__lane29_strm0_data_valid  ,

            // manager 53, lane 29, stream 1      
            input   wire                                        std__mgr53__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane29_strm1_data        ,
            output  wire                                        mgr53__std__lane29_strm1_data_valid  ,

            // manager 53, lane 30, stream 0      
            input   wire                                        std__mgr53__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane30_strm0_data        ,
            output  wire                                        mgr53__std__lane30_strm0_data_valid  ,

            // manager 53, lane 30, stream 1      
            input   wire                                        std__mgr53__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane30_strm1_data        ,
            output  wire                                        mgr53__std__lane30_strm1_data_valid  ,

            // manager 53, lane 31, stream 0      
            input   wire                                        std__mgr53__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane31_strm0_data        ,
            output  wire                                        mgr53__std__lane31_strm0_data_valid  ,

            // manager 53, lane 31, stream 1      
            input   wire                                        std__mgr53__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr53__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr53__std__lane31_strm1_data        ,
            output  wire                                        mgr53__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 54, lane 0, stream 0      
            input   wire                                        std__mgr54__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane0_strm0_data        ,
            output  wire                                        mgr54__std__lane0_strm0_data_valid  ,

            // manager 54, lane 0, stream 1      
            input   wire                                        std__mgr54__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane0_strm1_data        ,
            output  wire                                        mgr54__std__lane0_strm1_data_valid  ,

            // manager 54, lane 1, stream 0      
            input   wire                                        std__mgr54__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane1_strm0_data        ,
            output  wire                                        mgr54__std__lane1_strm0_data_valid  ,

            // manager 54, lane 1, stream 1      
            input   wire                                        std__mgr54__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane1_strm1_data        ,
            output  wire                                        mgr54__std__lane1_strm1_data_valid  ,

            // manager 54, lane 2, stream 0      
            input   wire                                        std__mgr54__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane2_strm0_data        ,
            output  wire                                        mgr54__std__lane2_strm0_data_valid  ,

            // manager 54, lane 2, stream 1      
            input   wire                                        std__mgr54__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane2_strm1_data        ,
            output  wire                                        mgr54__std__lane2_strm1_data_valid  ,

            // manager 54, lane 3, stream 0      
            input   wire                                        std__mgr54__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane3_strm0_data        ,
            output  wire                                        mgr54__std__lane3_strm0_data_valid  ,

            // manager 54, lane 3, stream 1      
            input   wire                                        std__mgr54__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane3_strm1_data        ,
            output  wire                                        mgr54__std__lane3_strm1_data_valid  ,

            // manager 54, lane 4, stream 0      
            input   wire                                        std__mgr54__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane4_strm0_data        ,
            output  wire                                        mgr54__std__lane4_strm0_data_valid  ,

            // manager 54, lane 4, stream 1      
            input   wire                                        std__mgr54__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane4_strm1_data        ,
            output  wire                                        mgr54__std__lane4_strm1_data_valid  ,

            // manager 54, lane 5, stream 0      
            input   wire                                        std__mgr54__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane5_strm0_data        ,
            output  wire                                        mgr54__std__lane5_strm0_data_valid  ,

            // manager 54, lane 5, stream 1      
            input   wire                                        std__mgr54__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane5_strm1_data        ,
            output  wire                                        mgr54__std__lane5_strm1_data_valid  ,

            // manager 54, lane 6, stream 0      
            input   wire                                        std__mgr54__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane6_strm0_data        ,
            output  wire                                        mgr54__std__lane6_strm0_data_valid  ,

            // manager 54, lane 6, stream 1      
            input   wire                                        std__mgr54__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane6_strm1_data        ,
            output  wire                                        mgr54__std__lane6_strm1_data_valid  ,

            // manager 54, lane 7, stream 0      
            input   wire                                        std__mgr54__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane7_strm0_data        ,
            output  wire                                        mgr54__std__lane7_strm0_data_valid  ,

            // manager 54, lane 7, stream 1      
            input   wire                                        std__mgr54__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane7_strm1_data        ,
            output  wire                                        mgr54__std__lane7_strm1_data_valid  ,

            // manager 54, lane 8, stream 0      
            input   wire                                        std__mgr54__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane8_strm0_data        ,
            output  wire                                        mgr54__std__lane8_strm0_data_valid  ,

            // manager 54, lane 8, stream 1      
            input   wire                                        std__mgr54__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane8_strm1_data        ,
            output  wire                                        mgr54__std__lane8_strm1_data_valid  ,

            // manager 54, lane 9, stream 0      
            input   wire                                        std__mgr54__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane9_strm0_data        ,
            output  wire                                        mgr54__std__lane9_strm0_data_valid  ,

            // manager 54, lane 9, stream 1      
            input   wire                                        std__mgr54__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane9_strm1_data        ,
            output  wire                                        mgr54__std__lane9_strm1_data_valid  ,

            // manager 54, lane 10, stream 0      
            input   wire                                        std__mgr54__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane10_strm0_data        ,
            output  wire                                        mgr54__std__lane10_strm0_data_valid  ,

            // manager 54, lane 10, stream 1      
            input   wire                                        std__mgr54__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane10_strm1_data        ,
            output  wire                                        mgr54__std__lane10_strm1_data_valid  ,

            // manager 54, lane 11, stream 0      
            input   wire                                        std__mgr54__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane11_strm0_data        ,
            output  wire                                        mgr54__std__lane11_strm0_data_valid  ,

            // manager 54, lane 11, stream 1      
            input   wire                                        std__mgr54__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane11_strm1_data        ,
            output  wire                                        mgr54__std__lane11_strm1_data_valid  ,

            // manager 54, lane 12, stream 0      
            input   wire                                        std__mgr54__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane12_strm0_data        ,
            output  wire                                        mgr54__std__lane12_strm0_data_valid  ,

            // manager 54, lane 12, stream 1      
            input   wire                                        std__mgr54__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane12_strm1_data        ,
            output  wire                                        mgr54__std__lane12_strm1_data_valid  ,

            // manager 54, lane 13, stream 0      
            input   wire                                        std__mgr54__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane13_strm0_data        ,
            output  wire                                        mgr54__std__lane13_strm0_data_valid  ,

            // manager 54, lane 13, stream 1      
            input   wire                                        std__mgr54__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane13_strm1_data        ,
            output  wire                                        mgr54__std__lane13_strm1_data_valid  ,

            // manager 54, lane 14, stream 0      
            input   wire                                        std__mgr54__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane14_strm0_data        ,
            output  wire                                        mgr54__std__lane14_strm0_data_valid  ,

            // manager 54, lane 14, stream 1      
            input   wire                                        std__mgr54__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane14_strm1_data        ,
            output  wire                                        mgr54__std__lane14_strm1_data_valid  ,

            // manager 54, lane 15, stream 0      
            input   wire                                        std__mgr54__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane15_strm0_data        ,
            output  wire                                        mgr54__std__lane15_strm0_data_valid  ,

            // manager 54, lane 15, stream 1      
            input   wire                                        std__mgr54__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane15_strm1_data        ,
            output  wire                                        mgr54__std__lane15_strm1_data_valid  ,

            // manager 54, lane 16, stream 0      
            input   wire                                        std__mgr54__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane16_strm0_data        ,
            output  wire                                        mgr54__std__lane16_strm0_data_valid  ,

            // manager 54, lane 16, stream 1      
            input   wire                                        std__mgr54__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane16_strm1_data        ,
            output  wire                                        mgr54__std__lane16_strm1_data_valid  ,

            // manager 54, lane 17, stream 0      
            input   wire                                        std__mgr54__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane17_strm0_data        ,
            output  wire                                        mgr54__std__lane17_strm0_data_valid  ,

            // manager 54, lane 17, stream 1      
            input   wire                                        std__mgr54__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane17_strm1_data        ,
            output  wire                                        mgr54__std__lane17_strm1_data_valid  ,

            // manager 54, lane 18, stream 0      
            input   wire                                        std__mgr54__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane18_strm0_data        ,
            output  wire                                        mgr54__std__lane18_strm0_data_valid  ,

            // manager 54, lane 18, stream 1      
            input   wire                                        std__mgr54__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane18_strm1_data        ,
            output  wire                                        mgr54__std__lane18_strm1_data_valid  ,

            // manager 54, lane 19, stream 0      
            input   wire                                        std__mgr54__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane19_strm0_data        ,
            output  wire                                        mgr54__std__lane19_strm0_data_valid  ,

            // manager 54, lane 19, stream 1      
            input   wire                                        std__mgr54__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane19_strm1_data        ,
            output  wire                                        mgr54__std__lane19_strm1_data_valid  ,

            // manager 54, lane 20, stream 0      
            input   wire                                        std__mgr54__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane20_strm0_data        ,
            output  wire                                        mgr54__std__lane20_strm0_data_valid  ,

            // manager 54, lane 20, stream 1      
            input   wire                                        std__mgr54__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane20_strm1_data        ,
            output  wire                                        mgr54__std__lane20_strm1_data_valid  ,

            // manager 54, lane 21, stream 0      
            input   wire                                        std__mgr54__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane21_strm0_data        ,
            output  wire                                        mgr54__std__lane21_strm0_data_valid  ,

            // manager 54, lane 21, stream 1      
            input   wire                                        std__mgr54__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane21_strm1_data        ,
            output  wire                                        mgr54__std__lane21_strm1_data_valid  ,

            // manager 54, lane 22, stream 0      
            input   wire                                        std__mgr54__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane22_strm0_data        ,
            output  wire                                        mgr54__std__lane22_strm0_data_valid  ,

            // manager 54, lane 22, stream 1      
            input   wire                                        std__mgr54__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane22_strm1_data        ,
            output  wire                                        mgr54__std__lane22_strm1_data_valid  ,

            // manager 54, lane 23, stream 0      
            input   wire                                        std__mgr54__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane23_strm0_data        ,
            output  wire                                        mgr54__std__lane23_strm0_data_valid  ,

            // manager 54, lane 23, stream 1      
            input   wire                                        std__mgr54__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane23_strm1_data        ,
            output  wire                                        mgr54__std__lane23_strm1_data_valid  ,

            // manager 54, lane 24, stream 0      
            input   wire                                        std__mgr54__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane24_strm0_data        ,
            output  wire                                        mgr54__std__lane24_strm0_data_valid  ,

            // manager 54, lane 24, stream 1      
            input   wire                                        std__mgr54__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane24_strm1_data        ,
            output  wire                                        mgr54__std__lane24_strm1_data_valid  ,

            // manager 54, lane 25, stream 0      
            input   wire                                        std__mgr54__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane25_strm0_data        ,
            output  wire                                        mgr54__std__lane25_strm0_data_valid  ,

            // manager 54, lane 25, stream 1      
            input   wire                                        std__mgr54__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane25_strm1_data        ,
            output  wire                                        mgr54__std__lane25_strm1_data_valid  ,

            // manager 54, lane 26, stream 0      
            input   wire                                        std__mgr54__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane26_strm0_data        ,
            output  wire                                        mgr54__std__lane26_strm0_data_valid  ,

            // manager 54, lane 26, stream 1      
            input   wire                                        std__mgr54__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane26_strm1_data        ,
            output  wire                                        mgr54__std__lane26_strm1_data_valid  ,

            // manager 54, lane 27, stream 0      
            input   wire                                        std__mgr54__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane27_strm0_data        ,
            output  wire                                        mgr54__std__lane27_strm0_data_valid  ,

            // manager 54, lane 27, stream 1      
            input   wire                                        std__mgr54__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane27_strm1_data        ,
            output  wire                                        mgr54__std__lane27_strm1_data_valid  ,

            // manager 54, lane 28, stream 0      
            input   wire                                        std__mgr54__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane28_strm0_data        ,
            output  wire                                        mgr54__std__lane28_strm0_data_valid  ,

            // manager 54, lane 28, stream 1      
            input   wire                                        std__mgr54__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane28_strm1_data        ,
            output  wire                                        mgr54__std__lane28_strm1_data_valid  ,

            // manager 54, lane 29, stream 0      
            input   wire                                        std__mgr54__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane29_strm0_data        ,
            output  wire                                        mgr54__std__lane29_strm0_data_valid  ,

            // manager 54, lane 29, stream 1      
            input   wire                                        std__mgr54__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane29_strm1_data        ,
            output  wire                                        mgr54__std__lane29_strm1_data_valid  ,

            // manager 54, lane 30, stream 0      
            input   wire                                        std__mgr54__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane30_strm0_data        ,
            output  wire                                        mgr54__std__lane30_strm0_data_valid  ,

            // manager 54, lane 30, stream 1      
            input   wire                                        std__mgr54__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane30_strm1_data        ,
            output  wire                                        mgr54__std__lane30_strm1_data_valid  ,

            // manager 54, lane 31, stream 0      
            input   wire                                        std__mgr54__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane31_strm0_data        ,
            output  wire                                        mgr54__std__lane31_strm0_data_valid  ,

            // manager 54, lane 31, stream 1      
            input   wire                                        std__mgr54__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr54__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr54__std__lane31_strm1_data        ,
            output  wire                                        mgr54__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 55, lane 0, stream 0      
            input   wire                                        std__mgr55__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane0_strm0_data        ,
            output  wire                                        mgr55__std__lane0_strm0_data_valid  ,

            // manager 55, lane 0, stream 1      
            input   wire                                        std__mgr55__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane0_strm1_data        ,
            output  wire                                        mgr55__std__lane0_strm1_data_valid  ,

            // manager 55, lane 1, stream 0      
            input   wire                                        std__mgr55__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane1_strm0_data        ,
            output  wire                                        mgr55__std__lane1_strm0_data_valid  ,

            // manager 55, lane 1, stream 1      
            input   wire                                        std__mgr55__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane1_strm1_data        ,
            output  wire                                        mgr55__std__lane1_strm1_data_valid  ,

            // manager 55, lane 2, stream 0      
            input   wire                                        std__mgr55__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane2_strm0_data        ,
            output  wire                                        mgr55__std__lane2_strm0_data_valid  ,

            // manager 55, lane 2, stream 1      
            input   wire                                        std__mgr55__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane2_strm1_data        ,
            output  wire                                        mgr55__std__lane2_strm1_data_valid  ,

            // manager 55, lane 3, stream 0      
            input   wire                                        std__mgr55__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane3_strm0_data        ,
            output  wire                                        mgr55__std__lane3_strm0_data_valid  ,

            // manager 55, lane 3, stream 1      
            input   wire                                        std__mgr55__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane3_strm1_data        ,
            output  wire                                        mgr55__std__lane3_strm1_data_valid  ,

            // manager 55, lane 4, stream 0      
            input   wire                                        std__mgr55__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane4_strm0_data        ,
            output  wire                                        mgr55__std__lane4_strm0_data_valid  ,

            // manager 55, lane 4, stream 1      
            input   wire                                        std__mgr55__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane4_strm1_data        ,
            output  wire                                        mgr55__std__lane4_strm1_data_valid  ,

            // manager 55, lane 5, stream 0      
            input   wire                                        std__mgr55__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane5_strm0_data        ,
            output  wire                                        mgr55__std__lane5_strm0_data_valid  ,

            // manager 55, lane 5, stream 1      
            input   wire                                        std__mgr55__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane5_strm1_data        ,
            output  wire                                        mgr55__std__lane5_strm1_data_valid  ,

            // manager 55, lane 6, stream 0      
            input   wire                                        std__mgr55__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane6_strm0_data        ,
            output  wire                                        mgr55__std__lane6_strm0_data_valid  ,

            // manager 55, lane 6, stream 1      
            input   wire                                        std__mgr55__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane6_strm1_data        ,
            output  wire                                        mgr55__std__lane6_strm1_data_valid  ,

            // manager 55, lane 7, stream 0      
            input   wire                                        std__mgr55__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane7_strm0_data        ,
            output  wire                                        mgr55__std__lane7_strm0_data_valid  ,

            // manager 55, lane 7, stream 1      
            input   wire                                        std__mgr55__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane7_strm1_data        ,
            output  wire                                        mgr55__std__lane7_strm1_data_valid  ,

            // manager 55, lane 8, stream 0      
            input   wire                                        std__mgr55__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane8_strm0_data        ,
            output  wire                                        mgr55__std__lane8_strm0_data_valid  ,

            // manager 55, lane 8, stream 1      
            input   wire                                        std__mgr55__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane8_strm1_data        ,
            output  wire                                        mgr55__std__lane8_strm1_data_valid  ,

            // manager 55, lane 9, stream 0      
            input   wire                                        std__mgr55__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane9_strm0_data        ,
            output  wire                                        mgr55__std__lane9_strm0_data_valid  ,

            // manager 55, lane 9, stream 1      
            input   wire                                        std__mgr55__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane9_strm1_data        ,
            output  wire                                        mgr55__std__lane9_strm1_data_valid  ,

            // manager 55, lane 10, stream 0      
            input   wire                                        std__mgr55__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane10_strm0_data        ,
            output  wire                                        mgr55__std__lane10_strm0_data_valid  ,

            // manager 55, lane 10, stream 1      
            input   wire                                        std__mgr55__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane10_strm1_data        ,
            output  wire                                        mgr55__std__lane10_strm1_data_valid  ,

            // manager 55, lane 11, stream 0      
            input   wire                                        std__mgr55__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane11_strm0_data        ,
            output  wire                                        mgr55__std__lane11_strm0_data_valid  ,

            // manager 55, lane 11, stream 1      
            input   wire                                        std__mgr55__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane11_strm1_data        ,
            output  wire                                        mgr55__std__lane11_strm1_data_valid  ,

            // manager 55, lane 12, stream 0      
            input   wire                                        std__mgr55__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane12_strm0_data        ,
            output  wire                                        mgr55__std__lane12_strm0_data_valid  ,

            // manager 55, lane 12, stream 1      
            input   wire                                        std__mgr55__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane12_strm1_data        ,
            output  wire                                        mgr55__std__lane12_strm1_data_valid  ,

            // manager 55, lane 13, stream 0      
            input   wire                                        std__mgr55__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane13_strm0_data        ,
            output  wire                                        mgr55__std__lane13_strm0_data_valid  ,

            // manager 55, lane 13, stream 1      
            input   wire                                        std__mgr55__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane13_strm1_data        ,
            output  wire                                        mgr55__std__lane13_strm1_data_valid  ,

            // manager 55, lane 14, stream 0      
            input   wire                                        std__mgr55__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane14_strm0_data        ,
            output  wire                                        mgr55__std__lane14_strm0_data_valid  ,

            // manager 55, lane 14, stream 1      
            input   wire                                        std__mgr55__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane14_strm1_data        ,
            output  wire                                        mgr55__std__lane14_strm1_data_valid  ,

            // manager 55, lane 15, stream 0      
            input   wire                                        std__mgr55__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane15_strm0_data        ,
            output  wire                                        mgr55__std__lane15_strm0_data_valid  ,

            // manager 55, lane 15, stream 1      
            input   wire                                        std__mgr55__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane15_strm1_data        ,
            output  wire                                        mgr55__std__lane15_strm1_data_valid  ,

            // manager 55, lane 16, stream 0      
            input   wire                                        std__mgr55__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane16_strm0_data        ,
            output  wire                                        mgr55__std__lane16_strm0_data_valid  ,

            // manager 55, lane 16, stream 1      
            input   wire                                        std__mgr55__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane16_strm1_data        ,
            output  wire                                        mgr55__std__lane16_strm1_data_valid  ,

            // manager 55, lane 17, stream 0      
            input   wire                                        std__mgr55__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane17_strm0_data        ,
            output  wire                                        mgr55__std__lane17_strm0_data_valid  ,

            // manager 55, lane 17, stream 1      
            input   wire                                        std__mgr55__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane17_strm1_data        ,
            output  wire                                        mgr55__std__lane17_strm1_data_valid  ,

            // manager 55, lane 18, stream 0      
            input   wire                                        std__mgr55__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane18_strm0_data        ,
            output  wire                                        mgr55__std__lane18_strm0_data_valid  ,

            // manager 55, lane 18, stream 1      
            input   wire                                        std__mgr55__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane18_strm1_data        ,
            output  wire                                        mgr55__std__lane18_strm1_data_valid  ,

            // manager 55, lane 19, stream 0      
            input   wire                                        std__mgr55__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane19_strm0_data        ,
            output  wire                                        mgr55__std__lane19_strm0_data_valid  ,

            // manager 55, lane 19, stream 1      
            input   wire                                        std__mgr55__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane19_strm1_data        ,
            output  wire                                        mgr55__std__lane19_strm1_data_valid  ,

            // manager 55, lane 20, stream 0      
            input   wire                                        std__mgr55__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane20_strm0_data        ,
            output  wire                                        mgr55__std__lane20_strm0_data_valid  ,

            // manager 55, lane 20, stream 1      
            input   wire                                        std__mgr55__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane20_strm1_data        ,
            output  wire                                        mgr55__std__lane20_strm1_data_valid  ,

            // manager 55, lane 21, stream 0      
            input   wire                                        std__mgr55__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane21_strm0_data        ,
            output  wire                                        mgr55__std__lane21_strm0_data_valid  ,

            // manager 55, lane 21, stream 1      
            input   wire                                        std__mgr55__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane21_strm1_data        ,
            output  wire                                        mgr55__std__lane21_strm1_data_valid  ,

            // manager 55, lane 22, stream 0      
            input   wire                                        std__mgr55__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane22_strm0_data        ,
            output  wire                                        mgr55__std__lane22_strm0_data_valid  ,

            // manager 55, lane 22, stream 1      
            input   wire                                        std__mgr55__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane22_strm1_data        ,
            output  wire                                        mgr55__std__lane22_strm1_data_valid  ,

            // manager 55, lane 23, stream 0      
            input   wire                                        std__mgr55__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane23_strm0_data        ,
            output  wire                                        mgr55__std__lane23_strm0_data_valid  ,

            // manager 55, lane 23, stream 1      
            input   wire                                        std__mgr55__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane23_strm1_data        ,
            output  wire                                        mgr55__std__lane23_strm1_data_valid  ,

            // manager 55, lane 24, stream 0      
            input   wire                                        std__mgr55__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane24_strm0_data        ,
            output  wire                                        mgr55__std__lane24_strm0_data_valid  ,

            // manager 55, lane 24, stream 1      
            input   wire                                        std__mgr55__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane24_strm1_data        ,
            output  wire                                        mgr55__std__lane24_strm1_data_valid  ,

            // manager 55, lane 25, stream 0      
            input   wire                                        std__mgr55__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane25_strm0_data        ,
            output  wire                                        mgr55__std__lane25_strm0_data_valid  ,

            // manager 55, lane 25, stream 1      
            input   wire                                        std__mgr55__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane25_strm1_data        ,
            output  wire                                        mgr55__std__lane25_strm1_data_valid  ,

            // manager 55, lane 26, stream 0      
            input   wire                                        std__mgr55__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane26_strm0_data        ,
            output  wire                                        mgr55__std__lane26_strm0_data_valid  ,

            // manager 55, lane 26, stream 1      
            input   wire                                        std__mgr55__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane26_strm1_data        ,
            output  wire                                        mgr55__std__lane26_strm1_data_valid  ,

            // manager 55, lane 27, stream 0      
            input   wire                                        std__mgr55__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane27_strm0_data        ,
            output  wire                                        mgr55__std__lane27_strm0_data_valid  ,

            // manager 55, lane 27, stream 1      
            input   wire                                        std__mgr55__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane27_strm1_data        ,
            output  wire                                        mgr55__std__lane27_strm1_data_valid  ,

            // manager 55, lane 28, stream 0      
            input   wire                                        std__mgr55__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane28_strm0_data        ,
            output  wire                                        mgr55__std__lane28_strm0_data_valid  ,

            // manager 55, lane 28, stream 1      
            input   wire                                        std__mgr55__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane28_strm1_data        ,
            output  wire                                        mgr55__std__lane28_strm1_data_valid  ,

            // manager 55, lane 29, stream 0      
            input   wire                                        std__mgr55__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane29_strm0_data        ,
            output  wire                                        mgr55__std__lane29_strm0_data_valid  ,

            // manager 55, lane 29, stream 1      
            input   wire                                        std__mgr55__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane29_strm1_data        ,
            output  wire                                        mgr55__std__lane29_strm1_data_valid  ,

            // manager 55, lane 30, stream 0      
            input   wire                                        std__mgr55__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane30_strm0_data        ,
            output  wire                                        mgr55__std__lane30_strm0_data_valid  ,

            // manager 55, lane 30, stream 1      
            input   wire                                        std__mgr55__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane30_strm1_data        ,
            output  wire                                        mgr55__std__lane30_strm1_data_valid  ,

            // manager 55, lane 31, stream 0      
            input   wire                                        std__mgr55__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane31_strm0_data        ,
            output  wire                                        mgr55__std__lane31_strm0_data_valid  ,

            // manager 55, lane 31, stream 1      
            input   wire                                        std__mgr55__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr55__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr55__std__lane31_strm1_data        ,
            output  wire                                        mgr55__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 56, lane 0, stream 0      
            input   wire                                        std__mgr56__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane0_strm0_data        ,
            output  wire                                        mgr56__std__lane0_strm0_data_valid  ,

            // manager 56, lane 0, stream 1      
            input   wire                                        std__mgr56__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane0_strm1_data        ,
            output  wire                                        mgr56__std__lane0_strm1_data_valid  ,

            // manager 56, lane 1, stream 0      
            input   wire                                        std__mgr56__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane1_strm0_data        ,
            output  wire                                        mgr56__std__lane1_strm0_data_valid  ,

            // manager 56, lane 1, stream 1      
            input   wire                                        std__mgr56__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane1_strm1_data        ,
            output  wire                                        mgr56__std__lane1_strm1_data_valid  ,

            // manager 56, lane 2, stream 0      
            input   wire                                        std__mgr56__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane2_strm0_data        ,
            output  wire                                        mgr56__std__lane2_strm0_data_valid  ,

            // manager 56, lane 2, stream 1      
            input   wire                                        std__mgr56__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane2_strm1_data        ,
            output  wire                                        mgr56__std__lane2_strm1_data_valid  ,

            // manager 56, lane 3, stream 0      
            input   wire                                        std__mgr56__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane3_strm0_data        ,
            output  wire                                        mgr56__std__lane3_strm0_data_valid  ,

            // manager 56, lane 3, stream 1      
            input   wire                                        std__mgr56__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane3_strm1_data        ,
            output  wire                                        mgr56__std__lane3_strm1_data_valid  ,

            // manager 56, lane 4, stream 0      
            input   wire                                        std__mgr56__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane4_strm0_data        ,
            output  wire                                        mgr56__std__lane4_strm0_data_valid  ,

            // manager 56, lane 4, stream 1      
            input   wire                                        std__mgr56__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane4_strm1_data        ,
            output  wire                                        mgr56__std__lane4_strm1_data_valid  ,

            // manager 56, lane 5, stream 0      
            input   wire                                        std__mgr56__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane5_strm0_data        ,
            output  wire                                        mgr56__std__lane5_strm0_data_valid  ,

            // manager 56, lane 5, stream 1      
            input   wire                                        std__mgr56__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane5_strm1_data        ,
            output  wire                                        mgr56__std__lane5_strm1_data_valid  ,

            // manager 56, lane 6, stream 0      
            input   wire                                        std__mgr56__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane6_strm0_data        ,
            output  wire                                        mgr56__std__lane6_strm0_data_valid  ,

            // manager 56, lane 6, stream 1      
            input   wire                                        std__mgr56__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane6_strm1_data        ,
            output  wire                                        mgr56__std__lane6_strm1_data_valid  ,

            // manager 56, lane 7, stream 0      
            input   wire                                        std__mgr56__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane7_strm0_data        ,
            output  wire                                        mgr56__std__lane7_strm0_data_valid  ,

            // manager 56, lane 7, stream 1      
            input   wire                                        std__mgr56__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane7_strm1_data        ,
            output  wire                                        mgr56__std__lane7_strm1_data_valid  ,

            // manager 56, lane 8, stream 0      
            input   wire                                        std__mgr56__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane8_strm0_data        ,
            output  wire                                        mgr56__std__lane8_strm0_data_valid  ,

            // manager 56, lane 8, stream 1      
            input   wire                                        std__mgr56__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane8_strm1_data        ,
            output  wire                                        mgr56__std__lane8_strm1_data_valid  ,

            // manager 56, lane 9, stream 0      
            input   wire                                        std__mgr56__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane9_strm0_data        ,
            output  wire                                        mgr56__std__lane9_strm0_data_valid  ,

            // manager 56, lane 9, stream 1      
            input   wire                                        std__mgr56__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane9_strm1_data        ,
            output  wire                                        mgr56__std__lane9_strm1_data_valid  ,

            // manager 56, lane 10, stream 0      
            input   wire                                        std__mgr56__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane10_strm0_data        ,
            output  wire                                        mgr56__std__lane10_strm0_data_valid  ,

            // manager 56, lane 10, stream 1      
            input   wire                                        std__mgr56__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane10_strm1_data        ,
            output  wire                                        mgr56__std__lane10_strm1_data_valid  ,

            // manager 56, lane 11, stream 0      
            input   wire                                        std__mgr56__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane11_strm0_data        ,
            output  wire                                        mgr56__std__lane11_strm0_data_valid  ,

            // manager 56, lane 11, stream 1      
            input   wire                                        std__mgr56__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane11_strm1_data        ,
            output  wire                                        mgr56__std__lane11_strm1_data_valid  ,

            // manager 56, lane 12, stream 0      
            input   wire                                        std__mgr56__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane12_strm0_data        ,
            output  wire                                        mgr56__std__lane12_strm0_data_valid  ,

            // manager 56, lane 12, stream 1      
            input   wire                                        std__mgr56__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane12_strm1_data        ,
            output  wire                                        mgr56__std__lane12_strm1_data_valid  ,

            // manager 56, lane 13, stream 0      
            input   wire                                        std__mgr56__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane13_strm0_data        ,
            output  wire                                        mgr56__std__lane13_strm0_data_valid  ,

            // manager 56, lane 13, stream 1      
            input   wire                                        std__mgr56__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane13_strm1_data        ,
            output  wire                                        mgr56__std__lane13_strm1_data_valid  ,

            // manager 56, lane 14, stream 0      
            input   wire                                        std__mgr56__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane14_strm0_data        ,
            output  wire                                        mgr56__std__lane14_strm0_data_valid  ,

            // manager 56, lane 14, stream 1      
            input   wire                                        std__mgr56__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane14_strm1_data        ,
            output  wire                                        mgr56__std__lane14_strm1_data_valid  ,

            // manager 56, lane 15, stream 0      
            input   wire                                        std__mgr56__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane15_strm0_data        ,
            output  wire                                        mgr56__std__lane15_strm0_data_valid  ,

            // manager 56, lane 15, stream 1      
            input   wire                                        std__mgr56__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane15_strm1_data        ,
            output  wire                                        mgr56__std__lane15_strm1_data_valid  ,

            // manager 56, lane 16, stream 0      
            input   wire                                        std__mgr56__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane16_strm0_data        ,
            output  wire                                        mgr56__std__lane16_strm0_data_valid  ,

            // manager 56, lane 16, stream 1      
            input   wire                                        std__mgr56__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane16_strm1_data        ,
            output  wire                                        mgr56__std__lane16_strm1_data_valid  ,

            // manager 56, lane 17, stream 0      
            input   wire                                        std__mgr56__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane17_strm0_data        ,
            output  wire                                        mgr56__std__lane17_strm0_data_valid  ,

            // manager 56, lane 17, stream 1      
            input   wire                                        std__mgr56__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane17_strm1_data        ,
            output  wire                                        mgr56__std__lane17_strm1_data_valid  ,

            // manager 56, lane 18, stream 0      
            input   wire                                        std__mgr56__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane18_strm0_data        ,
            output  wire                                        mgr56__std__lane18_strm0_data_valid  ,

            // manager 56, lane 18, stream 1      
            input   wire                                        std__mgr56__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane18_strm1_data        ,
            output  wire                                        mgr56__std__lane18_strm1_data_valid  ,

            // manager 56, lane 19, stream 0      
            input   wire                                        std__mgr56__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane19_strm0_data        ,
            output  wire                                        mgr56__std__lane19_strm0_data_valid  ,

            // manager 56, lane 19, stream 1      
            input   wire                                        std__mgr56__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane19_strm1_data        ,
            output  wire                                        mgr56__std__lane19_strm1_data_valid  ,

            // manager 56, lane 20, stream 0      
            input   wire                                        std__mgr56__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane20_strm0_data        ,
            output  wire                                        mgr56__std__lane20_strm0_data_valid  ,

            // manager 56, lane 20, stream 1      
            input   wire                                        std__mgr56__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane20_strm1_data        ,
            output  wire                                        mgr56__std__lane20_strm1_data_valid  ,

            // manager 56, lane 21, stream 0      
            input   wire                                        std__mgr56__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane21_strm0_data        ,
            output  wire                                        mgr56__std__lane21_strm0_data_valid  ,

            // manager 56, lane 21, stream 1      
            input   wire                                        std__mgr56__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane21_strm1_data        ,
            output  wire                                        mgr56__std__lane21_strm1_data_valid  ,

            // manager 56, lane 22, stream 0      
            input   wire                                        std__mgr56__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane22_strm0_data        ,
            output  wire                                        mgr56__std__lane22_strm0_data_valid  ,

            // manager 56, lane 22, stream 1      
            input   wire                                        std__mgr56__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane22_strm1_data        ,
            output  wire                                        mgr56__std__lane22_strm1_data_valid  ,

            // manager 56, lane 23, stream 0      
            input   wire                                        std__mgr56__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane23_strm0_data        ,
            output  wire                                        mgr56__std__lane23_strm0_data_valid  ,

            // manager 56, lane 23, stream 1      
            input   wire                                        std__mgr56__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane23_strm1_data        ,
            output  wire                                        mgr56__std__lane23_strm1_data_valid  ,

            // manager 56, lane 24, stream 0      
            input   wire                                        std__mgr56__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane24_strm0_data        ,
            output  wire                                        mgr56__std__lane24_strm0_data_valid  ,

            // manager 56, lane 24, stream 1      
            input   wire                                        std__mgr56__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane24_strm1_data        ,
            output  wire                                        mgr56__std__lane24_strm1_data_valid  ,

            // manager 56, lane 25, stream 0      
            input   wire                                        std__mgr56__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane25_strm0_data        ,
            output  wire                                        mgr56__std__lane25_strm0_data_valid  ,

            // manager 56, lane 25, stream 1      
            input   wire                                        std__mgr56__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane25_strm1_data        ,
            output  wire                                        mgr56__std__lane25_strm1_data_valid  ,

            // manager 56, lane 26, stream 0      
            input   wire                                        std__mgr56__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane26_strm0_data        ,
            output  wire                                        mgr56__std__lane26_strm0_data_valid  ,

            // manager 56, lane 26, stream 1      
            input   wire                                        std__mgr56__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane26_strm1_data        ,
            output  wire                                        mgr56__std__lane26_strm1_data_valid  ,

            // manager 56, lane 27, stream 0      
            input   wire                                        std__mgr56__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane27_strm0_data        ,
            output  wire                                        mgr56__std__lane27_strm0_data_valid  ,

            // manager 56, lane 27, stream 1      
            input   wire                                        std__mgr56__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane27_strm1_data        ,
            output  wire                                        mgr56__std__lane27_strm1_data_valid  ,

            // manager 56, lane 28, stream 0      
            input   wire                                        std__mgr56__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane28_strm0_data        ,
            output  wire                                        mgr56__std__lane28_strm0_data_valid  ,

            // manager 56, lane 28, stream 1      
            input   wire                                        std__mgr56__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane28_strm1_data        ,
            output  wire                                        mgr56__std__lane28_strm1_data_valid  ,

            // manager 56, lane 29, stream 0      
            input   wire                                        std__mgr56__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane29_strm0_data        ,
            output  wire                                        mgr56__std__lane29_strm0_data_valid  ,

            // manager 56, lane 29, stream 1      
            input   wire                                        std__mgr56__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane29_strm1_data        ,
            output  wire                                        mgr56__std__lane29_strm1_data_valid  ,

            // manager 56, lane 30, stream 0      
            input   wire                                        std__mgr56__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane30_strm0_data        ,
            output  wire                                        mgr56__std__lane30_strm0_data_valid  ,

            // manager 56, lane 30, stream 1      
            input   wire                                        std__mgr56__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane30_strm1_data        ,
            output  wire                                        mgr56__std__lane30_strm1_data_valid  ,

            // manager 56, lane 31, stream 0      
            input   wire                                        std__mgr56__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane31_strm0_data        ,
            output  wire                                        mgr56__std__lane31_strm0_data_valid  ,

            // manager 56, lane 31, stream 1      
            input   wire                                        std__mgr56__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr56__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr56__std__lane31_strm1_data        ,
            output  wire                                        mgr56__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 57, lane 0, stream 0      
            input   wire                                        std__mgr57__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane0_strm0_data        ,
            output  wire                                        mgr57__std__lane0_strm0_data_valid  ,

            // manager 57, lane 0, stream 1      
            input   wire                                        std__mgr57__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane0_strm1_data        ,
            output  wire                                        mgr57__std__lane0_strm1_data_valid  ,

            // manager 57, lane 1, stream 0      
            input   wire                                        std__mgr57__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane1_strm0_data        ,
            output  wire                                        mgr57__std__lane1_strm0_data_valid  ,

            // manager 57, lane 1, stream 1      
            input   wire                                        std__mgr57__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane1_strm1_data        ,
            output  wire                                        mgr57__std__lane1_strm1_data_valid  ,

            // manager 57, lane 2, stream 0      
            input   wire                                        std__mgr57__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane2_strm0_data        ,
            output  wire                                        mgr57__std__lane2_strm0_data_valid  ,

            // manager 57, lane 2, stream 1      
            input   wire                                        std__mgr57__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane2_strm1_data        ,
            output  wire                                        mgr57__std__lane2_strm1_data_valid  ,

            // manager 57, lane 3, stream 0      
            input   wire                                        std__mgr57__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane3_strm0_data        ,
            output  wire                                        mgr57__std__lane3_strm0_data_valid  ,

            // manager 57, lane 3, stream 1      
            input   wire                                        std__mgr57__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane3_strm1_data        ,
            output  wire                                        mgr57__std__lane3_strm1_data_valid  ,

            // manager 57, lane 4, stream 0      
            input   wire                                        std__mgr57__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane4_strm0_data        ,
            output  wire                                        mgr57__std__lane4_strm0_data_valid  ,

            // manager 57, lane 4, stream 1      
            input   wire                                        std__mgr57__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane4_strm1_data        ,
            output  wire                                        mgr57__std__lane4_strm1_data_valid  ,

            // manager 57, lane 5, stream 0      
            input   wire                                        std__mgr57__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane5_strm0_data        ,
            output  wire                                        mgr57__std__lane5_strm0_data_valid  ,

            // manager 57, lane 5, stream 1      
            input   wire                                        std__mgr57__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane5_strm1_data        ,
            output  wire                                        mgr57__std__lane5_strm1_data_valid  ,

            // manager 57, lane 6, stream 0      
            input   wire                                        std__mgr57__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane6_strm0_data        ,
            output  wire                                        mgr57__std__lane6_strm0_data_valid  ,

            // manager 57, lane 6, stream 1      
            input   wire                                        std__mgr57__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane6_strm1_data        ,
            output  wire                                        mgr57__std__lane6_strm1_data_valid  ,

            // manager 57, lane 7, stream 0      
            input   wire                                        std__mgr57__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane7_strm0_data        ,
            output  wire                                        mgr57__std__lane7_strm0_data_valid  ,

            // manager 57, lane 7, stream 1      
            input   wire                                        std__mgr57__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane7_strm1_data        ,
            output  wire                                        mgr57__std__lane7_strm1_data_valid  ,

            // manager 57, lane 8, stream 0      
            input   wire                                        std__mgr57__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane8_strm0_data        ,
            output  wire                                        mgr57__std__lane8_strm0_data_valid  ,

            // manager 57, lane 8, stream 1      
            input   wire                                        std__mgr57__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane8_strm1_data        ,
            output  wire                                        mgr57__std__lane8_strm1_data_valid  ,

            // manager 57, lane 9, stream 0      
            input   wire                                        std__mgr57__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane9_strm0_data        ,
            output  wire                                        mgr57__std__lane9_strm0_data_valid  ,

            // manager 57, lane 9, stream 1      
            input   wire                                        std__mgr57__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane9_strm1_data        ,
            output  wire                                        mgr57__std__lane9_strm1_data_valid  ,

            // manager 57, lane 10, stream 0      
            input   wire                                        std__mgr57__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane10_strm0_data        ,
            output  wire                                        mgr57__std__lane10_strm0_data_valid  ,

            // manager 57, lane 10, stream 1      
            input   wire                                        std__mgr57__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane10_strm1_data        ,
            output  wire                                        mgr57__std__lane10_strm1_data_valid  ,

            // manager 57, lane 11, stream 0      
            input   wire                                        std__mgr57__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane11_strm0_data        ,
            output  wire                                        mgr57__std__lane11_strm0_data_valid  ,

            // manager 57, lane 11, stream 1      
            input   wire                                        std__mgr57__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane11_strm1_data        ,
            output  wire                                        mgr57__std__lane11_strm1_data_valid  ,

            // manager 57, lane 12, stream 0      
            input   wire                                        std__mgr57__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane12_strm0_data        ,
            output  wire                                        mgr57__std__lane12_strm0_data_valid  ,

            // manager 57, lane 12, stream 1      
            input   wire                                        std__mgr57__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane12_strm1_data        ,
            output  wire                                        mgr57__std__lane12_strm1_data_valid  ,

            // manager 57, lane 13, stream 0      
            input   wire                                        std__mgr57__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane13_strm0_data        ,
            output  wire                                        mgr57__std__lane13_strm0_data_valid  ,

            // manager 57, lane 13, stream 1      
            input   wire                                        std__mgr57__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane13_strm1_data        ,
            output  wire                                        mgr57__std__lane13_strm1_data_valid  ,

            // manager 57, lane 14, stream 0      
            input   wire                                        std__mgr57__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane14_strm0_data        ,
            output  wire                                        mgr57__std__lane14_strm0_data_valid  ,

            // manager 57, lane 14, stream 1      
            input   wire                                        std__mgr57__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane14_strm1_data        ,
            output  wire                                        mgr57__std__lane14_strm1_data_valid  ,

            // manager 57, lane 15, stream 0      
            input   wire                                        std__mgr57__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane15_strm0_data        ,
            output  wire                                        mgr57__std__lane15_strm0_data_valid  ,

            // manager 57, lane 15, stream 1      
            input   wire                                        std__mgr57__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane15_strm1_data        ,
            output  wire                                        mgr57__std__lane15_strm1_data_valid  ,

            // manager 57, lane 16, stream 0      
            input   wire                                        std__mgr57__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane16_strm0_data        ,
            output  wire                                        mgr57__std__lane16_strm0_data_valid  ,

            // manager 57, lane 16, stream 1      
            input   wire                                        std__mgr57__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane16_strm1_data        ,
            output  wire                                        mgr57__std__lane16_strm1_data_valid  ,

            // manager 57, lane 17, stream 0      
            input   wire                                        std__mgr57__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane17_strm0_data        ,
            output  wire                                        mgr57__std__lane17_strm0_data_valid  ,

            // manager 57, lane 17, stream 1      
            input   wire                                        std__mgr57__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane17_strm1_data        ,
            output  wire                                        mgr57__std__lane17_strm1_data_valid  ,

            // manager 57, lane 18, stream 0      
            input   wire                                        std__mgr57__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane18_strm0_data        ,
            output  wire                                        mgr57__std__lane18_strm0_data_valid  ,

            // manager 57, lane 18, stream 1      
            input   wire                                        std__mgr57__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane18_strm1_data        ,
            output  wire                                        mgr57__std__lane18_strm1_data_valid  ,

            // manager 57, lane 19, stream 0      
            input   wire                                        std__mgr57__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane19_strm0_data        ,
            output  wire                                        mgr57__std__lane19_strm0_data_valid  ,

            // manager 57, lane 19, stream 1      
            input   wire                                        std__mgr57__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane19_strm1_data        ,
            output  wire                                        mgr57__std__lane19_strm1_data_valid  ,

            // manager 57, lane 20, stream 0      
            input   wire                                        std__mgr57__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane20_strm0_data        ,
            output  wire                                        mgr57__std__lane20_strm0_data_valid  ,

            // manager 57, lane 20, stream 1      
            input   wire                                        std__mgr57__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane20_strm1_data        ,
            output  wire                                        mgr57__std__lane20_strm1_data_valid  ,

            // manager 57, lane 21, stream 0      
            input   wire                                        std__mgr57__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane21_strm0_data        ,
            output  wire                                        mgr57__std__lane21_strm0_data_valid  ,

            // manager 57, lane 21, stream 1      
            input   wire                                        std__mgr57__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane21_strm1_data        ,
            output  wire                                        mgr57__std__lane21_strm1_data_valid  ,

            // manager 57, lane 22, stream 0      
            input   wire                                        std__mgr57__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane22_strm0_data        ,
            output  wire                                        mgr57__std__lane22_strm0_data_valid  ,

            // manager 57, lane 22, stream 1      
            input   wire                                        std__mgr57__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane22_strm1_data        ,
            output  wire                                        mgr57__std__lane22_strm1_data_valid  ,

            // manager 57, lane 23, stream 0      
            input   wire                                        std__mgr57__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane23_strm0_data        ,
            output  wire                                        mgr57__std__lane23_strm0_data_valid  ,

            // manager 57, lane 23, stream 1      
            input   wire                                        std__mgr57__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane23_strm1_data        ,
            output  wire                                        mgr57__std__lane23_strm1_data_valid  ,

            // manager 57, lane 24, stream 0      
            input   wire                                        std__mgr57__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane24_strm0_data        ,
            output  wire                                        mgr57__std__lane24_strm0_data_valid  ,

            // manager 57, lane 24, stream 1      
            input   wire                                        std__mgr57__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane24_strm1_data        ,
            output  wire                                        mgr57__std__lane24_strm1_data_valid  ,

            // manager 57, lane 25, stream 0      
            input   wire                                        std__mgr57__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane25_strm0_data        ,
            output  wire                                        mgr57__std__lane25_strm0_data_valid  ,

            // manager 57, lane 25, stream 1      
            input   wire                                        std__mgr57__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane25_strm1_data        ,
            output  wire                                        mgr57__std__lane25_strm1_data_valid  ,

            // manager 57, lane 26, stream 0      
            input   wire                                        std__mgr57__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane26_strm0_data        ,
            output  wire                                        mgr57__std__lane26_strm0_data_valid  ,

            // manager 57, lane 26, stream 1      
            input   wire                                        std__mgr57__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane26_strm1_data        ,
            output  wire                                        mgr57__std__lane26_strm1_data_valid  ,

            // manager 57, lane 27, stream 0      
            input   wire                                        std__mgr57__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane27_strm0_data        ,
            output  wire                                        mgr57__std__lane27_strm0_data_valid  ,

            // manager 57, lane 27, stream 1      
            input   wire                                        std__mgr57__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane27_strm1_data        ,
            output  wire                                        mgr57__std__lane27_strm1_data_valid  ,

            // manager 57, lane 28, stream 0      
            input   wire                                        std__mgr57__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane28_strm0_data        ,
            output  wire                                        mgr57__std__lane28_strm0_data_valid  ,

            // manager 57, lane 28, stream 1      
            input   wire                                        std__mgr57__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane28_strm1_data        ,
            output  wire                                        mgr57__std__lane28_strm1_data_valid  ,

            // manager 57, lane 29, stream 0      
            input   wire                                        std__mgr57__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane29_strm0_data        ,
            output  wire                                        mgr57__std__lane29_strm0_data_valid  ,

            // manager 57, lane 29, stream 1      
            input   wire                                        std__mgr57__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane29_strm1_data        ,
            output  wire                                        mgr57__std__lane29_strm1_data_valid  ,

            // manager 57, lane 30, stream 0      
            input   wire                                        std__mgr57__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane30_strm0_data        ,
            output  wire                                        mgr57__std__lane30_strm0_data_valid  ,

            // manager 57, lane 30, stream 1      
            input   wire                                        std__mgr57__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane30_strm1_data        ,
            output  wire                                        mgr57__std__lane30_strm1_data_valid  ,

            // manager 57, lane 31, stream 0      
            input   wire                                        std__mgr57__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane31_strm0_data        ,
            output  wire                                        mgr57__std__lane31_strm0_data_valid  ,

            // manager 57, lane 31, stream 1      
            input   wire                                        std__mgr57__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr57__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr57__std__lane31_strm1_data        ,
            output  wire                                        mgr57__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 58, lane 0, stream 0      
            input   wire                                        std__mgr58__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane0_strm0_data        ,
            output  wire                                        mgr58__std__lane0_strm0_data_valid  ,

            // manager 58, lane 0, stream 1      
            input   wire                                        std__mgr58__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane0_strm1_data        ,
            output  wire                                        mgr58__std__lane0_strm1_data_valid  ,

            // manager 58, lane 1, stream 0      
            input   wire                                        std__mgr58__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane1_strm0_data        ,
            output  wire                                        mgr58__std__lane1_strm0_data_valid  ,

            // manager 58, lane 1, stream 1      
            input   wire                                        std__mgr58__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane1_strm1_data        ,
            output  wire                                        mgr58__std__lane1_strm1_data_valid  ,

            // manager 58, lane 2, stream 0      
            input   wire                                        std__mgr58__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane2_strm0_data        ,
            output  wire                                        mgr58__std__lane2_strm0_data_valid  ,

            // manager 58, lane 2, stream 1      
            input   wire                                        std__mgr58__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane2_strm1_data        ,
            output  wire                                        mgr58__std__lane2_strm1_data_valid  ,

            // manager 58, lane 3, stream 0      
            input   wire                                        std__mgr58__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane3_strm0_data        ,
            output  wire                                        mgr58__std__lane3_strm0_data_valid  ,

            // manager 58, lane 3, stream 1      
            input   wire                                        std__mgr58__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane3_strm1_data        ,
            output  wire                                        mgr58__std__lane3_strm1_data_valid  ,

            // manager 58, lane 4, stream 0      
            input   wire                                        std__mgr58__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane4_strm0_data        ,
            output  wire                                        mgr58__std__lane4_strm0_data_valid  ,

            // manager 58, lane 4, stream 1      
            input   wire                                        std__mgr58__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane4_strm1_data        ,
            output  wire                                        mgr58__std__lane4_strm1_data_valid  ,

            // manager 58, lane 5, stream 0      
            input   wire                                        std__mgr58__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane5_strm0_data        ,
            output  wire                                        mgr58__std__lane5_strm0_data_valid  ,

            // manager 58, lane 5, stream 1      
            input   wire                                        std__mgr58__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane5_strm1_data        ,
            output  wire                                        mgr58__std__lane5_strm1_data_valid  ,

            // manager 58, lane 6, stream 0      
            input   wire                                        std__mgr58__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane6_strm0_data        ,
            output  wire                                        mgr58__std__lane6_strm0_data_valid  ,

            // manager 58, lane 6, stream 1      
            input   wire                                        std__mgr58__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane6_strm1_data        ,
            output  wire                                        mgr58__std__lane6_strm1_data_valid  ,

            // manager 58, lane 7, stream 0      
            input   wire                                        std__mgr58__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane7_strm0_data        ,
            output  wire                                        mgr58__std__lane7_strm0_data_valid  ,

            // manager 58, lane 7, stream 1      
            input   wire                                        std__mgr58__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane7_strm1_data        ,
            output  wire                                        mgr58__std__lane7_strm1_data_valid  ,

            // manager 58, lane 8, stream 0      
            input   wire                                        std__mgr58__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane8_strm0_data        ,
            output  wire                                        mgr58__std__lane8_strm0_data_valid  ,

            // manager 58, lane 8, stream 1      
            input   wire                                        std__mgr58__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane8_strm1_data        ,
            output  wire                                        mgr58__std__lane8_strm1_data_valid  ,

            // manager 58, lane 9, stream 0      
            input   wire                                        std__mgr58__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane9_strm0_data        ,
            output  wire                                        mgr58__std__lane9_strm0_data_valid  ,

            // manager 58, lane 9, stream 1      
            input   wire                                        std__mgr58__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane9_strm1_data        ,
            output  wire                                        mgr58__std__lane9_strm1_data_valid  ,

            // manager 58, lane 10, stream 0      
            input   wire                                        std__mgr58__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane10_strm0_data        ,
            output  wire                                        mgr58__std__lane10_strm0_data_valid  ,

            // manager 58, lane 10, stream 1      
            input   wire                                        std__mgr58__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane10_strm1_data        ,
            output  wire                                        mgr58__std__lane10_strm1_data_valid  ,

            // manager 58, lane 11, stream 0      
            input   wire                                        std__mgr58__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane11_strm0_data        ,
            output  wire                                        mgr58__std__lane11_strm0_data_valid  ,

            // manager 58, lane 11, stream 1      
            input   wire                                        std__mgr58__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane11_strm1_data        ,
            output  wire                                        mgr58__std__lane11_strm1_data_valid  ,

            // manager 58, lane 12, stream 0      
            input   wire                                        std__mgr58__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane12_strm0_data        ,
            output  wire                                        mgr58__std__lane12_strm0_data_valid  ,

            // manager 58, lane 12, stream 1      
            input   wire                                        std__mgr58__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane12_strm1_data        ,
            output  wire                                        mgr58__std__lane12_strm1_data_valid  ,

            // manager 58, lane 13, stream 0      
            input   wire                                        std__mgr58__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane13_strm0_data        ,
            output  wire                                        mgr58__std__lane13_strm0_data_valid  ,

            // manager 58, lane 13, stream 1      
            input   wire                                        std__mgr58__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane13_strm1_data        ,
            output  wire                                        mgr58__std__lane13_strm1_data_valid  ,

            // manager 58, lane 14, stream 0      
            input   wire                                        std__mgr58__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane14_strm0_data        ,
            output  wire                                        mgr58__std__lane14_strm0_data_valid  ,

            // manager 58, lane 14, stream 1      
            input   wire                                        std__mgr58__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane14_strm1_data        ,
            output  wire                                        mgr58__std__lane14_strm1_data_valid  ,

            // manager 58, lane 15, stream 0      
            input   wire                                        std__mgr58__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane15_strm0_data        ,
            output  wire                                        mgr58__std__lane15_strm0_data_valid  ,

            // manager 58, lane 15, stream 1      
            input   wire                                        std__mgr58__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane15_strm1_data        ,
            output  wire                                        mgr58__std__lane15_strm1_data_valid  ,

            // manager 58, lane 16, stream 0      
            input   wire                                        std__mgr58__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane16_strm0_data        ,
            output  wire                                        mgr58__std__lane16_strm0_data_valid  ,

            // manager 58, lane 16, stream 1      
            input   wire                                        std__mgr58__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane16_strm1_data        ,
            output  wire                                        mgr58__std__lane16_strm1_data_valid  ,

            // manager 58, lane 17, stream 0      
            input   wire                                        std__mgr58__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane17_strm0_data        ,
            output  wire                                        mgr58__std__lane17_strm0_data_valid  ,

            // manager 58, lane 17, stream 1      
            input   wire                                        std__mgr58__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane17_strm1_data        ,
            output  wire                                        mgr58__std__lane17_strm1_data_valid  ,

            // manager 58, lane 18, stream 0      
            input   wire                                        std__mgr58__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane18_strm0_data        ,
            output  wire                                        mgr58__std__lane18_strm0_data_valid  ,

            // manager 58, lane 18, stream 1      
            input   wire                                        std__mgr58__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane18_strm1_data        ,
            output  wire                                        mgr58__std__lane18_strm1_data_valid  ,

            // manager 58, lane 19, stream 0      
            input   wire                                        std__mgr58__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane19_strm0_data        ,
            output  wire                                        mgr58__std__lane19_strm0_data_valid  ,

            // manager 58, lane 19, stream 1      
            input   wire                                        std__mgr58__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane19_strm1_data        ,
            output  wire                                        mgr58__std__lane19_strm1_data_valid  ,

            // manager 58, lane 20, stream 0      
            input   wire                                        std__mgr58__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane20_strm0_data        ,
            output  wire                                        mgr58__std__lane20_strm0_data_valid  ,

            // manager 58, lane 20, stream 1      
            input   wire                                        std__mgr58__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane20_strm1_data        ,
            output  wire                                        mgr58__std__lane20_strm1_data_valid  ,

            // manager 58, lane 21, stream 0      
            input   wire                                        std__mgr58__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane21_strm0_data        ,
            output  wire                                        mgr58__std__lane21_strm0_data_valid  ,

            // manager 58, lane 21, stream 1      
            input   wire                                        std__mgr58__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane21_strm1_data        ,
            output  wire                                        mgr58__std__lane21_strm1_data_valid  ,

            // manager 58, lane 22, stream 0      
            input   wire                                        std__mgr58__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane22_strm0_data        ,
            output  wire                                        mgr58__std__lane22_strm0_data_valid  ,

            // manager 58, lane 22, stream 1      
            input   wire                                        std__mgr58__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane22_strm1_data        ,
            output  wire                                        mgr58__std__lane22_strm1_data_valid  ,

            // manager 58, lane 23, stream 0      
            input   wire                                        std__mgr58__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane23_strm0_data        ,
            output  wire                                        mgr58__std__lane23_strm0_data_valid  ,

            // manager 58, lane 23, stream 1      
            input   wire                                        std__mgr58__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane23_strm1_data        ,
            output  wire                                        mgr58__std__lane23_strm1_data_valid  ,

            // manager 58, lane 24, stream 0      
            input   wire                                        std__mgr58__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane24_strm0_data        ,
            output  wire                                        mgr58__std__lane24_strm0_data_valid  ,

            // manager 58, lane 24, stream 1      
            input   wire                                        std__mgr58__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane24_strm1_data        ,
            output  wire                                        mgr58__std__lane24_strm1_data_valid  ,

            // manager 58, lane 25, stream 0      
            input   wire                                        std__mgr58__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane25_strm0_data        ,
            output  wire                                        mgr58__std__lane25_strm0_data_valid  ,

            // manager 58, lane 25, stream 1      
            input   wire                                        std__mgr58__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane25_strm1_data        ,
            output  wire                                        mgr58__std__lane25_strm1_data_valid  ,

            // manager 58, lane 26, stream 0      
            input   wire                                        std__mgr58__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane26_strm0_data        ,
            output  wire                                        mgr58__std__lane26_strm0_data_valid  ,

            // manager 58, lane 26, stream 1      
            input   wire                                        std__mgr58__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane26_strm1_data        ,
            output  wire                                        mgr58__std__lane26_strm1_data_valid  ,

            // manager 58, lane 27, stream 0      
            input   wire                                        std__mgr58__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane27_strm0_data        ,
            output  wire                                        mgr58__std__lane27_strm0_data_valid  ,

            // manager 58, lane 27, stream 1      
            input   wire                                        std__mgr58__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane27_strm1_data        ,
            output  wire                                        mgr58__std__lane27_strm1_data_valid  ,

            // manager 58, lane 28, stream 0      
            input   wire                                        std__mgr58__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane28_strm0_data        ,
            output  wire                                        mgr58__std__lane28_strm0_data_valid  ,

            // manager 58, lane 28, stream 1      
            input   wire                                        std__mgr58__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane28_strm1_data        ,
            output  wire                                        mgr58__std__lane28_strm1_data_valid  ,

            // manager 58, lane 29, stream 0      
            input   wire                                        std__mgr58__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane29_strm0_data        ,
            output  wire                                        mgr58__std__lane29_strm0_data_valid  ,

            // manager 58, lane 29, stream 1      
            input   wire                                        std__mgr58__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane29_strm1_data        ,
            output  wire                                        mgr58__std__lane29_strm1_data_valid  ,

            // manager 58, lane 30, stream 0      
            input   wire                                        std__mgr58__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane30_strm0_data        ,
            output  wire                                        mgr58__std__lane30_strm0_data_valid  ,

            // manager 58, lane 30, stream 1      
            input   wire                                        std__mgr58__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane30_strm1_data        ,
            output  wire                                        mgr58__std__lane30_strm1_data_valid  ,

            // manager 58, lane 31, stream 0      
            input   wire                                        std__mgr58__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane31_strm0_data        ,
            output  wire                                        mgr58__std__lane31_strm0_data_valid  ,

            // manager 58, lane 31, stream 1      
            input   wire                                        std__mgr58__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr58__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr58__std__lane31_strm1_data        ,
            output  wire                                        mgr58__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 59, lane 0, stream 0      
            input   wire                                        std__mgr59__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane0_strm0_data        ,
            output  wire                                        mgr59__std__lane0_strm0_data_valid  ,

            // manager 59, lane 0, stream 1      
            input   wire                                        std__mgr59__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane0_strm1_data        ,
            output  wire                                        mgr59__std__lane0_strm1_data_valid  ,

            // manager 59, lane 1, stream 0      
            input   wire                                        std__mgr59__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane1_strm0_data        ,
            output  wire                                        mgr59__std__lane1_strm0_data_valid  ,

            // manager 59, lane 1, stream 1      
            input   wire                                        std__mgr59__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane1_strm1_data        ,
            output  wire                                        mgr59__std__lane1_strm1_data_valid  ,

            // manager 59, lane 2, stream 0      
            input   wire                                        std__mgr59__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane2_strm0_data        ,
            output  wire                                        mgr59__std__lane2_strm0_data_valid  ,

            // manager 59, lane 2, stream 1      
            input   wire                                        std__mgr59__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane2_strm1_data        ,
            output  wire                                        mgr59__std__lane2_strm1_data_valid  ,

            // manager 59, lane 3, stream 0      
            input   wire                                        std__mgr59__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane3_strm0_data        ,
            output  wire                                        mgr59__std__lane3_strm0_data_valid  ,

            // manager 59, lane 3, stream 1      
            input   wire                                        std__mgr59__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane3_strm1_data        ,
            output  wire                                        mgr59__std__lane3_strm1_data_valid  ,

            // manager 59, lane 4, stream 0      
            input   wire                                        std__mgr59__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane4_strm0_data        ,
            output  wire                                        mgr59__std__lane4_strm0_data_valid  ,

            // manager 59, lane 4, stream 1      
            input   wire                                        std__mgr59__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane4_strm1_data        ,
            output  wire                                        mgr59__std__lane4_strm1_data_valid  ,

            // manager 59, lane 5, stream 0      
            input   wire                                        std__mgr59__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane5_strm0_data        ,
            output  wire                                        mgr59__std__lane5_strm0_data_valid  ,

            // manager 59, lane 5, stream 1      
            input   wire                                        std__mgr59__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane5_strm1_data        ,
            output  wire                                        mgr59__std__lane5_strm1_data_valid  ,

            // manager 59, lane 6, stream 0      
            input   wire                                        std__mgr59__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane6_strm0_data        ,
            output  wire                                        mgr59__std__lane6_strm0_data_valid  ,

            // manager 59, lane 6, stream 1      
            input   wire                                        std__mgr59__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane6_strm1_data        ,
            output  wire                                        mgr59__std__lane6_strm1_data_valid  ,

            // manager 59, lane 7, stream 0      
            input   wire                                        std__mgr59__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane7_strm0_data        ,
            output  wire                                        mgr59__std__lane7_strm0_data_valid  ,

            // manager 59, lane 7, stream 1      
            input   wire                                        std__mgr59__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane7_strm1_data        ,
            output  wire                                        mgr59__std__lane7_strm1_data_valid  ,

            // manager 59, lane 8, stream 0      
            input   wire                                        std__mgr59__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane8_strm0_data        ,
            output  wire                                        mgr59__std__lane8_strm0_data_valid  ,

            // manager 59, lane 8, stream 1      
            input   wire                                        std__mgr59__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane8_strm1_data        ,
            output  wire                                        mgr59__std__lane8_strm1_data_valid  ,

            // manager 59, lane 9, stream 0      
            input   wire                                        std__mgr59__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane9_strm0_data        ,
            output  wire                                        mgr59__std__lane9_strm0_data_valid  ,

            // manager 59, lane 9, stream 1      
            input   wire                                        std__mgr59__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane9_strm1_data        ,
            output  wire                                        mgr59__std__lane9_strm1_data_valid  ,

            // manager 59, lane 10, stream 0      
            input   wire                                        std__mgr59__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane10_strm0_data        ,
            output  wire                                        mgr59__std__lane10_strm0_data_valid  ,

            // manager 59, lane 10, stream 1      
            input   wire                                        std__mgr59__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane10_strm1_data        ,
            output  wire                                        mgr59__std__lane10_strm1_data_valid  ,

            // manager 59, lane 11, stream 0      
            input   wire                                        std__mgr59__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane11_strm0_data        ,
            output  wire                                        mgr59__std__lane11_strm0_data_valid  ,

            // manager 59, lane 11, stream 1      
            input   wire                                        std__mgr59__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane11_strm1_data        ,
            output  wire                                        mgr59__std__lane11_strm1_data_valid  ,

            // manager 59, lane 12, stream 0      
            input   wire                                        std__mgr59__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane12_strm0_data        ,
            output  wire                                        mgr59__std__lane12_strm0_data_valid  ,

            // manager 59, lane 12, stream 1      
            input   wire                                        std__mgr59__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane12_strm1_data        ,
            output  wire                                        mgr59__std__lane12_strm1_data_valid  ,

            // manager 59, lane 13, stream 0      
            input   wire                                        std__mgr59__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane13_strm0_data        ,
            output  wire                                        mgr59__std__lane13_strm0_data_valid  ,

            // manager 59, lane 13, stream 1      
            input   wire                                        std__mgr59__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane13_strm1_data        ,
            output  wire                                        mgr59__std__lane13_strm1_data_valid  ,

            // manager 59, lane 14, stream 0      
            input   wire                                        std__mgr59__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane14_strm0_data        ,
            output  wire                                        mgr59__std__lane14_strm0_data_valid  ,

            // manager 59, lane 14, stream 1      
            input   wire                                        std__mgr59__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane14_strm1_data        ,
            output  wire                                        mgr59__std__lane14_strm1_data_valid  ,

            // manager 59, lane 15, stream 0      
            input   wire                                        std__mgr59__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane15_strm0_data        ,
            output  wire                                        mgr59__std__lane15_strm0_data_valid  ,

            // manager 59, lane 15, stream 1      
            input   wire                                        std__mgr59__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane15_strm1_data        ,
            output  wire                                        mgr59__std__lane15_strm1_data_valid  ,

            // manager 59, lane 16, stream 0      
            input   wire                                        std__mgr59__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane16_strm0_data        ,
            output  wire                                        mgr59__std__lane16_strm0_data_valid  ,

            // manager 59, lane 16, stream 1      
            input   wire                                        std__mgr59__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane16_strm1_data        ,
            output  wire                                        mgr59__std__lane16_strm1_data_valid  ,

            // manager 59, lane 17, stream 0      
            input   wire                                        std__mgr59__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane17_strm0_data        ,
            output  wire                                        mgr59__std__lane17_strm0_data_valid  ,

            // manager 59, lane 17, stream 1      
            input   wire                                        std__mgr59__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane17_strm1_data        ,
            output  wire                                        mgr59__std__lane17_strm1_data_valid  ,

            // manager 59, lane 18, stream 0      
            input   wire                                        std__mgr59__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane18_strm0_data        ,
            output  wire                                        mgr59__std__lane18_strm0_data_valid  ,

            // manager 59, lane 18, stream 1      
            input   wire                                        std__mgr59__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane18_strm1_data        ,
            output  wire                                        mgr59__std__lane18_strm1_data_valid  ,

            // manager 59, lane 19, stream 0      
            input   wire                                        std__mgr59__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane19_strm0_data        ,
            output  wire                                        mgr59__std__lane19_strm0_data_valid  ,

            // manager 59, lane 19, stream 1      
            input   wire                                        std__mgr59__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane19_strm1_data        ,
            output  wire                                        mgr59__std__lane19_strm1_data_valid  ,

            // manager 59, lane 20, stream 0      
            input   wire                                        std__mgr59__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane20_strm0_data        ,
            output  wire                                        mgr59__std__lane20_strm0_data_valid  ,

            // manager 59, lane 20, stream 1      
            input   wire                                        std__mgr59__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane20_strm1_data        ,
            output  wire                                        mgr59__std__lane20_strm1_data_valid  ,

            // manager 59, lane 21, stream 0      
            input   wire                                        std__mgr59__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane21_strm0_data        ,
            output  wire                                        mgr59__std__lane21_strm0_data_valid  ,

            // manager 59, lane 21, stream 1      
            input   wire                                        std__mgr59__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane21_strm1_data        ,
            output  wire                                        mgr59__std__lane21_strm1_data_valid  ,

            // manager 59, lane 22, stream 0      
            input   wire                                        std__mgr59__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane22_strm0_data        ,
            output  wire                                        mgr59__std__lane22_strm0_data_valid  ,

            // manager 59, lane 22, stream 1      
            input   wire                                        std__mgr59__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane22_strm1_data        ,
            output  wire                                        mgr59__std__lane22_strm1_data_valid  ,

            // manager 59, lane 23, stream 0      
            input   wire                                        std__mgr59__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane23_strm0_data        ,
            output  wire                                        mgr59__std__lane23_strm0_data_valid  ,

            // manager 59, lane 23, stream 1      
            input   wire                                        std__mgr59__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane23_strm1_data        ,
            output  wire                                        mgr59__std__lane23_strm1_data_valid  ,

            // manager 59, lane 24, stream 0      
            input   wire                                        std__mgr59__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane24_strm0_data        ,
            output  wire                                        mgr59__std__lane24_strm0_data_valid  ,

            // manager 59, lane 24, stream 1      
            input   wire                                        std__mgr59__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane24_strm1_data        ,
            output  wire                                        mgr59__std__lane24_strm1_data_valid  ,

            // manager 59, lane 25, stream 0      
            input   wire                                        std__mgr59__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane25_strm0_data        ,
            output  wire                                        mgr59__std__lane25_strm0_data_valid  ,

            // manager 59, lane 25, stream 1      
            input   wire                                        std__mgr59__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane25_strm1_data        ,
            output  wire                                        mgr59__std__lane25_strm1_data_valid  ,

            // manager 59, lane 26, stream 0      
            input   wire                                        std__mgr59__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane26_strm0_data        ,
            output  wire                                        mgr59__std__lane26_strm0_data_valid  ,

            // manager 59, lane 26, stream 1      
            input   wire                                        std__mgr59__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane26_strm1_data        ,
            output  wire                                        mgr59__std__lane26_strm1_data_valid  ,

            // manager 59, lane 27, stream 0      
            input   wire                                        std__mgr59__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane27_strm0_data        ,
            output  wire                                        mgr59__std__lane27_strm0_data_valid  ,

            // manager 59, lane 27, stream 1      
            input   wire                                        std__mgr59__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane27_strm1_data        ,
            output  wire                                        mgr59__std__lane27_strm1_data_valid  ,

            // manager 59, lane 28, stream 0      
            input   wire                                        std__mgr59__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane28_strm0_data        ,
            output  wire                                        mgr59__std__lane28_strm0_data_valid  ,

            // manager 59, lane 28, stream 1      
            input   wire                                        std__mgr59__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane28_strm1_data        ,
            output  wire                                        mgr59__std__lane28_strm1_data_valid  ,

            // manager 59, lane 29, stream 0      
            input   wire                                        std__mgr59__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane29_strm0_data        ,
            output  wire                                        mgr59__std__lane29_strm0_data_valid  ,

            // manager 59, lane 29, stream 1      
            input   wire                                        std__mgr59__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane29_strm1_data        ,
            output  wire                                        mgr59__std__lane29_strm1_data_valid  ,

            // manager 59, lane 30, stream 0      
            input   wire                                        std__mgr59__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane30_strm0_data        ,
            output  wire                                        mgr59__std__lane30_strm0_data_valid  ,

            // manager 59, lane 30, stream 1      
            input   wire                                        std__mgr59__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane30_strm1_data        ,
            output  wire                                        mgr59__std__lane30_strm1_data_valid  ,

            // manager 59, lane 31, stream 0      
            input   wire                                        std__mgr59__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane31_strm0_data        ,
            output  wire                                        mgr59__std__lane31_strm0_data_valid  ,

            // manager 59, lane 31, stream 1      
            input   wire                                        std__mgr59__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr59__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr59__std__lane31_strm1_data        ,
            output  wire                                        mgr59__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 60, lane 0, stream 0      
            input   wire                                        std__mgr60__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane0_strm0_data        ,
            output  wire                                        mgr60__std__lane0_strm0_data_valid  ,

            // manager 60, lane 0, stream 1      
            input   wire                                        std__mgr60__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane0_strm1_data        ,
            output  wire                                        mgr60__std__lane0_strm1_data_valid  ,

            // manager 60, lane 1, stream 0      
            input   wire                                        std__mgr60__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane1_strm0_data        ,
            output  wire                                        mgr60__std__lane1_strm0_data_valid  ,

            // manager 60, lane 1, stream 1      
            input   wire                                        std__mgr60__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane1_strm1_data        ,
            output  wire                                        mgr60__std__lane1_strm1_data_valid  ,

            // manager 60, lane 2, stream 0      
            input   wire                                        std__mgr60__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane2_strm0_data        ,
            output  wire                                        mgr60__std__lane2_strm0_data_valid  ,

            // manager 60, lane 2, stream 1      
            input   wire                                        std__mgr60__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane2_strm1_data        ,
            output  wire                                        mgr60__std__lane2_strm1_data_valid  ,

            // manager 60, lane 3, stream 0      
            input   wire                                        std__mgr60__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane3_strm0_data        ,
            output  wire                                        mgr60__std__lane3_strm0_data_valid  ,

            // manager 60, lane 3, stream 1      
            input   wire                                        std__mgr60__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane3_strm1_data        ,
            output  wire                                        mgr60__std__lane3_strm1_data_valid  ,

            // manager 60, lane 4, stream 0      
            input   wire                                        std__mgr60__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane4_strm0_data        ,
            output  wire                                        mgr60__std__lane4_strm0_data_valid  ,

            // manager 60, lane 4, stream 1      
            input   wire                                        std__mgr60__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane4_strm1_data        ,
            output  wire                                        mgr60__std__lane4_strm1_data_valid  ,

            // manager 60, lane 5, stream 0      
            input   wire                                        std__mgr60__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane5_strm0_data        ,
            output  wire                                        mgr60__std__lane5_strm0_data_valid  ,

            // manager 60, lane 5, stream 1      
            input   wire                                        std__mgr60__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane5_strm1_data        ,
            output  wire                                        mgr60__std__lane5_strm1_data_valid  ,

            // manager 60, lane 6, stream 0      
            input   wire                                        std__mgr60__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane6_strm0_data        ,
            output  wire                                        mgr60__std__lane6_strm0_data_valid  ,

            // manager 60, lane 6, stream 1      
            input   wire                                        std__mgr60__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane6_strm1_data        ,
            output  wire                                        mgr60__std__lane6_strm1_data_valid  ,

            // manager 60, lane 7, stream 0      
            input   wire                                        std__mgr60__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane7_strm0_data        ,
            output  wire                                        mgr60__std__lane7_strm0_data_valid  ,

            // manager 60, lane 7, stream 1      
            input   wire                                        std__mgr60__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane7_strm1_data        ,
            output  wire                                        mgr60__std__lane7_strm1_data_valid  ,

            // manager 60, lane 8, stream 0      
            input   wire                                        std__mgr60__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane8_strm0_data        ,
            output  wire                                        mgr60__std__lane8_strm0_data_valid  ,

            // manager 60, lane 8, stream 1      
            input   wire                                        std__mgr60__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane8_strm1_data        ,
            output  wire                                        mgr60__std__lane8_strm1_data_valid  ,

            // manager 60, lane 9, stream 0      
            input   wire                                        std__mgr60__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane9_strm0_data        ,
            output  wire                                        mgr60__std__lane9_strm0_data_valid  ,

            // manager 60, lane 9, stream 1      
            input   wire                                        std__mgr60__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane9_strm1_data        ,
            output  wire                                        mgr60__std__lane9_strm1_data_valid  ,

            // manager 60, lane 10, stream 0      
            input   wire                                        std__mgr60__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane10_strm0_data        ,
            output  wire                                        mgr60__std__lane10_strm0_data_valid  ,

            // manager 60, lane 10, stream 1      
            input   wire                                        std__mgr60__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane10_strm1_data        ,
            output  wire                                        mgr60__std__lane10_strm1_data_valid  ,

            // manager 60, lane 11, stream 0      
            input   wire                                        std__mgr60__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane11_strm0_data        ,
            output  wire                                        mgr60__std__lane11_strm0_data_valid  ,

            // manager 60, lane 11, stream 1      
            input   wire                                        std__mgr60__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane11_strm1_data        ,
            output  wire                                        mgr60__std__lane11_strm1_data_valid  ,

            // manager 60, lane 12, stream 0      
            input   wire                                        std__mgr60__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane12_strm0_data        ,
            output  wire                                        mgr60__std__lane12_strm0_data_valid  ,

            // manager 60, lane 12, stream 1      
            input   wire                                        std__mgr60__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane12_strm1_data        ,
            output  wire                                        mgr60__std__lane12_strm1_data_valid  ,

            // manager 60, lane 13, stream 0      
            input   wire                                        std__mgr60__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane13_strm0_data        ,
            output  wire                                        mgr60__std__lane13_strm0_data_valid  ,

            // manager 60, lane 13, stream 1      
            input   wire                                        std__mgr60__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane13_strm1_data        ,
            output  wire                                        mgr60__std__lane13_strm1_data_valid  ,

            // manager 60, lane 14, stream 0      
            input   wire                                        std__mgr60__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane14_strm0_data        ,
            output  wire                                        mgr60__std__lane14_strm0_data_valid  ,

            // manager 60, lane 14, stream 1      
            input   wire                                        std__mgr60__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane14_strm1_data        ,
            output  wire                                        mgr60__std__lane14_strm1_data_valid  ,

            // manager 60, lane 15, stream 0      
            input   wire                                        std__mgr60__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane15_strm0_data        ,
            output  wire                                        mgr60__std__lane15_strm0_data_valid  ,

            // manager 60, lane 15, stream 1      
            input   wire                                        std__mgr60__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane15_strm1_data        ,
            output  wire                                        mgr60__std__lane15_strm1_data_valid  ,

            // manager 60, lane 16, stream 0      
            input   wire                                        std__mgr60__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane16_strm0_data        ,
            output  wire                                        mgr60__std__lane16_strm0_data_valid  ,

            // manager 60, lane 16, stream 1      
            input   wire                                        std__mgr60__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane16_strm1_data        ,
            output  wire                                        mgr60__std__lane16_strm1_data_valid  ,

            // manager 60, lane 17, stream 0      
            input   wire                                        std__mgr60__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane17_strm0_data        ,
            output  wire                                        mgr60__std__lane17_strm0_data_valid  ,

            // manager 60, lane 17, stream 1      
            input   wire                                        std__mgr60__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane17_strm1_data        ,
            output  wire                                        mgr60__std__lane17_strm1_data_valid  ,

            // manager 60, lane 18, stream 0      
            input   wire                                        std__mgr60__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane18_strm0_data        ,
            output  wire                                        mgr60__std__lane18_strm0_data_valid  ,

            // manager 60, lane 18, stream 1      
            input   wire                                        std__mgr60__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane18_strm1_data        ,
            output  wire                                        mgr60__std__lane18_strm1_data_valid  ,

            // manager 60, lane 19, stream 0      
            input   wire                                        std__mgr60__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane19_strm0_data        ,
            output  wire                                        mgr60__std__lane19_strm0_data_valid  ,

            // manager 60, lane 19, stream 1      
            input   wire                                        std__mgr60__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane19_strm1_data        ,
            output  wire                                        mgr60__std__lane19_strm1_data_valid  ,

            // manager 60, lane 20, stream 0      
            input   wire                                        std__mgr60__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane20_strm0_data        ,
            output  wire                                        mgr60__std__lane20_strm0_data_valid  ,

            // manager 60, lane 20, stream 1      
            input   wire                                        std__mgr60__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane20_strm1_data        ,
            output  wire                                        mgr60__std__lane20_strm1_data_valid  ,

            // manager 60, lane 21, stream 0      
            input   wire                                        std__mgr60__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane21_strm0_data        ,
            output  wire                                        mgr60__std__lane21_strm0_data_valid  ,

            // manager 60, lane 21, stream 1      
            input   wire                                        std__mgr60__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane21_strm1_data        ,
            output  wire                                        mgr60__std__lane21_strm1_data_valid  ,

            // manager 60, lane 22, stream 0      
            input   wire                                        std__mgr60__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane22_strm0_data        ,
            output  wire                                        mgr60__std__lane22_strm0_data_valid  ,

            // manager 60, lane 22, stream 1      
            input   wire                                        std__mgr60__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane22_strm1_data        ,
            output  wire                                        mgr60__std__lane22_strm1_data_valid  ,

            // manager 60, lane 23, stream 0      
            input   wire                                        std__mgr60__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane23_strm0_data        ,
            output  wire                                        mgr60__std__lane23_strm0_data_valid  ,

            // manager 60, lane 23, stream 1      
            input   wire                                        std__mgr60__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane23_strm1_data        ,
            output  wire                                        mgr60__std__lane23_strm1_data_valid  ,

            // manager 60, lane 24, stream 0      
            input   wire                                        std__mgr60__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane24_strm0_data        ,
            output  wire                                        mgr60__std__lane24_strm0_data_valid  ,

            // manager 60, lane 24, stream 1      
            input   wire                                        std__mgr60__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane24_strm1_data        ,
            output  wire                                        mgr60__std__lane24_strm1_data_valid  ,

            // manager 60, lane 25, stream 0      
            input   wire                                        std__mgr60__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane25_strm0_data        ,
            output  wire                                        mgr60__std__lane25_strm0_data_valid  ,

            // manager 60, lane 25, stream 1      
            input   wire                                        std__mgr60__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane25_strm1_data        ,
            output  wire                                        mgr60__std__lane25_strm1_data_valid  ,

            // manager 60, lane 26, stream 0      
            input   wire                                        std__mgr60__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane26_strm0_data        ,
            output  wire                                        mgr60__std__lane26_strm0_data_valid  ,

            // manager 60, lane 26, stream 1      
            input   wire                                        std__mgr60__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane26_strm1_data        ,
            output  wire                                        mgr60__std__lane26_strm1_data_valid  ,

            // manager 60, lane 27, stream 0      
            input   wire                                        std__mgr60__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane27_strm0_data        ,
            output  wire                                        mgr60__std__lane27_strm0_data_valid  ,

            // manager 60, lane 27, stream 1      
            input   wire                                        std__mgr60__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane27_strm1_data        ,
            output  wire                                        mgr60__std__lane27_strm1_data_valid  ,

            // manager 60, lane 28, stream 0      
            input   wire                                        std__mgr60__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane28_strm0_data        ,
            output  wire                                        mgr60__std__lane28_strm0_data_valid  ,

            // manager 60, lane 28, stream 1      
            input   wire                                        std__mgr60__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane28_strm1_data        ,
            output  wire                                        mgr60__std__lane28_strm1_data_valid  ,

            // manager 60, lane 29, stream 0      
            input   wire                                        std__mgr60__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane29_strm0_data        ,
            output  wire                                        mgr60__std__lane29_strm0_data_valid  ,

            // manager 60, lane 29, stream 1      
            input   wire                                        std__mgr60__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane29_strm1_data        ,
            output  wire                                        mgr60__std__lane29_strm1_data_valid  ,

            // manager 60, lane 30, stream 0      
            input   wire                                        std__mgr60__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane30_strm0_data        ,
            output  wire                                        mgr60__std__lane30_strm0_data_valid  ,

            // manager 60, lane 30, stream 1      
            input   wire                                        std__mgr60__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane30_strm1_data        ,
            output  wire                                        mgr60__std__lane30_strm1_data_valid  ,

            // manager 60, lane 31, stream 0      
            input   wire                                        std__mgr60__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane31_strm0_data        ,
            output  wire                                        mgr60__std__lane31_strm0_data_valid  ,

            // manager 60, lane 31, stream 1      
            input   wire                                        std__mgr60__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr60__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr60__std__lane31_strm1_data        ,
            output  wire                                        mgr60__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 61, lane 0, stream 0      
            input   wire                                        std__mgr61__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane0_strm0_data        ,
            output  wire                                        mgr61__std__lane0_strm0_data_valid  ,

            // manager 61, lane 0, stream 1      
            input   wire                                        std__mgr61__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane0_strm1_data        ,
            output  wire                                        mgr61__std__lane0_strm1_data_valid  ,

            // manager 61, lane 1, stream 0      
            input   wire                                        std__mgr61__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane1_strm0_data        ,
            output  wire                                        mgr61__std__lane1_strm0_data_valid  ,

            // manager 61, lane 1, stream 1      
            input   wire                                        std__mgr61__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane1_strm1_data        ,
            output  wire                                        mgr61__std__lane1_strm1_data_valid  ,

            // manager 61, lane 2, stream 0      
            input   wire                                        std__mgr61__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane2_strm0_data        ,
            output  wire                                        mgr61__std__lane2_strm0_data_valid  ,

            // manager 61, lane 2, stream 1      
            input   wire                                        std__mgr61__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane2_strm1_data        ,
            output  wire                                        mgr61__std__lane2_strm1_data_valid  ,

            // manager 61, lane 3, stream 0      
            input   wire                                        std__mgr61__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane3_strm0_data        ,
            output  wire                                        mgr61__std__lane3_strm0_data_valid  ,

            // manager 61, lane 3, stream 1      
            input   wire                                        std__mgr61__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane3_strm1_data        ,
            output  wire                                        mgr61__std__lane3_strm1_data_valid  ,

            // manager 61, lane 4, stream 0      
            input   wire                                        std__mgr61__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane4_strm0_data        ,
            output  wire                                        mgr61__std__lane4_strm0_data_valid  ,

            // manager 61, lane 4, stream 1      
            input   wire                                        std__mgr61__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane4_strm1_data        ,
            output  wire                                        mgr61__std__lane4_strm1_data_valid  ,

            // manager 61, lane 5, stream 0      
            input   wire                                        std__mgr61__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane5_strm0_data        ,
            output  wire                                        mgr61__std__lane5_strm0_data_valid  ,

            // manager 61, lane 5, stream 1      
            input   wire                                        std__mgr61__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane5_strm1_data        ,
            output  wire                                        mgr61__std__lane5_strm1_data_valid  ,

            // manager 61, lane 6, stream 0      
            input   wire                                        std__mgr61__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane6_strm0_data        ,
            output  wire                                        mgr61__std__lane6_strm0_data_valid  ,

            // manager 61, lane 6, stream 1      
            input   wire                                        std__mgr61__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane6_strm1_data        ,
            output  wire                                        mgr61__std__lane6_strm1_data_valid  ,

            // manager 61, lane 7, stream 0      
            input   wire                                        std__mgr61__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane7_strm0_data        ,
            output  wire                                        mgr61__std__lane7_strm0_data_valid  ,

            // manager 61, lane 7, stream 1      
            input   wire                                        std__mgr61__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane7_strm1_data        ,
            output  wire                                        mgr61__std__lane7_strm1_data_valid  ,

            // manager 61, lane 8, stream 0      
            input   wire                                        std__mgr61__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane8_strm0_data        ,
            output  wire                                        mgr61__std__lane8_strm0_data_valid  ,

            // manager 61, lane 8, stream 1      
            input   wire                                        std__mgr61__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane8_strm1_data        ,
            output  wire                                        mgr61__std__lane8_strm1_data_valid  ,

            // manager 61, lane 9, stream 0      
            input   wire                                        std__mgr61__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane9_strm0_data        ,
            output  wire                                        mgr61__std__lane9_strm0_data_valid  ,

            // manager 61, lane 9, stream 1      
            input   wire                                        std__mgr61__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane9_strm1_data        ,
            output  wire                                        mgr61__std__lane9_strm1_data_valid  ,

            // manager 61, lane 10, stream 0      
            input   wire                                        std__mgr61__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane10_strm0_data        ,
            output  wire                                        mgr61__std__lane10_strm0_data_valid  ,

            // manager 61, lane 10, stream 1      
            input   wire                                        std__mgr61__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane10_strm1_data        ,
            output  wire                                        mgr61__std__lane10_strm1_data_valid  ,

            // manager 61, lane 11, stream 0      
            input   wire                                        std__mgr61__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane11_strm0_data        ,
            output  wire                                        mgr61__std__lane11_strm0_data_valid  ,

            // manager 61, lane 11, stream 1      
            input   wire                                        std__mgr61__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane11_strm1_data        ,
            output  wire                                        mgr61__std__lane11_strm1_data_valid  ,

            // manager 61, lane 12, stream 0      
            input   wire                                        std__mgr61__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane12_strm0_data        ,
            output  wire                                        mgr61__std__lane12_strm0_data_valid  ,

            // manager 61, lane 12, stream 1      
            input   wire                                        std__mgr61__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane12_strm1_data        ,
            output  wire                                        mgr61__std__lane12_strm1_data_valid  ,

            // manager 61, lane 13, stream 0      
            input   wire                                        std__mgr61__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane13_strm0_data        ,
            output  wire                                        mgr61__std__lane13_strm0_data_valid  ,

            // manager 61, lane 13, stream 1      
            input   wire                                        std__mgr61__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane13_strm1_data        ,
            output  wire                                        mgr61__std__lane13_strm1_data_valid  ,

            // manager 61, lane 14, stream 0      
            input   wire                                        std__mgr61__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane14_strm0_data        ,
            output  wire                                        mgr61__std__lane14_strm0_data_valid  ,

            // manager 61, lane 14, stream 1      
            input   wire                                        std__mgr61__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane14_strm1_data        ,
            output  wire                                        mgr61__std__lane14_strm1_data_valid  ,

            // manager 61, lane 15, stream 0      
            input   wire                                        std__mgr61__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane15_strm0_data        ,
            output  wire                                        mgr61__std__lane15_strm0_data_valid  ,

            // manager 61, lane 15, stream 1      
            input   wire                                        std__mgr61__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane15_strm1_data        ,
            output  wire                                        mgr61__std__lane15_strm1_data_valid  ,

            // manager 61, lane 16, stream 0      
            input   wire                                        std__mgr61__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane16_strm0_data        ,
            output  wire                                        mgr61__std__lane16_strm0_data_valid  ,

            // manager 61, lane 16, stream 1      
            input   wire                                        std__mgr61__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane16_strm1_data        ,
            output  wire                                        mgr61__std__lane16_strm1_data_valid  ,

            // manager 61, lane 17, stream 0      
            input   wire                                        std__mgr61__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane17_strm0_data        ,
            output  wire                                        mgr61__std__lane17_strm0_data_valid  ,

            // manager 61, lane 17, stream 1      
            input   wire                                        std__mgr61__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane17_strm1_data        ,
            output  wire                                        mgr61__std__lane17_strm1_data_valid  ,

            // manager 61, lane 18, stream 0      
            input   wire                                        std__mgr61__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane18_strm0_data        ,
            output  wire                                        mgr61__std__lane18_strm0_data_valid  ,

            // manager 61, lane 18, stream 1      
            input   wire                                        std__mgr61__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane18_strm1_data        ,
            output  wire                                        mgr61__std__lane18_strm1_data_valid  ,

            // manager 61, lane 19, stream 0      
            input   wire                                        std__mgr61__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane19_strm0_data        ,
            output  wire                                        mgr61__std__lane19_strm0_data_valid  ,

            // manager 61, lane 19, stream 1      
            input   wire                                        std__mgr61__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane19_strm1_data        ,
            output  wire                                        mgr61__std__lane19_strm1_data_valid  ,

            // manager 61, lane 20, stream 0      
            input   wire                                        std__mgr61__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane20_strm0_data        ,
            output  wire                                        mgr61__std__lane20_strm0_data_valid  ,

            // manager 61, lane 20, stream 1      
            input   wire                                        std__mgr61__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane20_strm1_data        ,
            output  wire                                        mgr61__std__lane20_strm1_data_valid  ,

            // manager 61, lane 21, stream 0      
            input   wire                                        std__mgr61__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane21_strm0_data        ,
            output  wire                                        mgr61__std__lane21_strm0_data_valid  ,

            // manager 61, lane 21, stream 1      
            input   wire                                        std__mgr61__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane21_strm1_data        ,
            output  wire                                        mgr61__std__lane21_strm1_data_valid  ,

            // manager 61, lane 22, stream 0      
            input   wire                                        std__mgr61__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane22_strm0_data        ,
            output  wire                                        mgr61__std__lane22_strm0_data_valid  ,

            // manager 61, lane 22, stream 1      
            input   wire                                        std__mgr61__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane22_strm1_data        ,
            output  wire                                        mgr61__std__lane22_strm1_data_valid  ,

            // manager 61, lane 23, stream 0      
            input   wire                                        std__mgr61__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane23_strm0_data        ,
            output  wire                                        mgr61__std__lane23_strm0_data_valid  ,

            // manager 61, lane 23, stream 1      
            input   wire                                        std__mgr61__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane23_strm1_data        ,
            output  wire                                        mgr61__std__lane23_strm1_data_valid  ,

            // manager 61, lane 24, stream 0      
            input   wire                                        std__mgr61__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane24_strm0_data        ,
            output  wire                                        mgr61__std__lane24_strm0_data_valid  ,

            // manager 61, lane 24, stream 1      
            input   wire                                        std__mgr61__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane24_strm1_data        ,
            output  wire                                        mgr61__std__lane24_strm1_data_valid  ,

            // manager 61, lane 25, stream 0      
            input   wire                                        std__mgr61__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane25_strm0_data        ,
            output  wire                                        mgr61__std__lane25_strm0_data_valid  ,

            // manager 61, lane 25, stream 1      
            input   wire                                        std__mgr61__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane25_strm1_data        ,
            output  wire                                        mgr61__std__lane25_strm1_data_valid  ,

            // manager 61, lane 26, stream 0      
            input   wire                                        std__mgr61__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane26_strm0_data        ,
            output  wire                                        mgr61__std__lane26_strm0_data_valid  ,

            // manager 61, lane 26, stream 1      
            input   wire                                        std__mgr61__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane26_strm1_data        ,
            output  wire                                        mgr61__std__lane26_strm1_data_valid  ,

            // manager 61, lane 27, stream 0      
            input   wire                                        std__mgr61__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane27_strm0_data        ,
            output  wire                                        mgr61__std__lane27_strm0_data_valid  ,

            // manager 61, lane 27, stream 1      
            input   wire                                        std__mgr61__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane27_strm1_data        ,
            output  wire                                        mgr61__std__lane27_strm1_data_valid  ,

            // manager 61, lane 28, stream 0      
            input   wire                                        std__mgr61__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane28_strm0_data        ,
            output  wire                                        mgr61__std__lane28_strm0_data_valid  ,

            // manager 61, lane 28, stream 1      
            input   wire                                        std__mgr61__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane28_strm1_data        ,
            output  wire                                        mgr61__std__lane28_strm1_data_valid  ,

            // manager 61, lane 29, stream 0      
            input   wire                                        std__mgr61__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane29_strm0_data        ,
            output  wire                                        mgr61__std__lane29_strm0_data_valid  ,

            // manager 61, lane 29, stream 1      
            input   wire                                        std__mgr61__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane29_strm1_data        ,
            output  wire                                        mgr61__std__lane29_strm1_data_valid  ,

            // manager 61, lane 30, stream 0      
            input   wire                                        std__mgr61__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane30_strm0_data        ,
            output  wire                                        mgr61__std__lane30_strm0_data_valid  ,

            // manager 61, lane 30, stream 1      
            input   wire                                        std__mgr61__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane30_strm1_data        ,
            output  wire                                        mgr61__std__lane30_strm1_data_valid  ,

            // manager 61, lane 31, stream 0      
            input   wire                                        std__mgr61__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane31_strm0_data        ,
            output  wire                                        mgr61__std__lane31_strm0_data_valid  ,

            // manager 61, lane 31, stream 1      
            input   wire                                        std__mgr61__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr61__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr61__std__lane31_strm1_data        ,
            output  wire                                        mgr61__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 62, lane 0, stream 0      
            input   wire                                        std__mgr62__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane0_strm0_data        ,
            output  wire                                        mgr62__std__lane0_strm0_data_valid  ,

            // manager 62, lane 0, stream 1      
            input   wire                                        std__mgr62__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane0_strm1_data        ,
            output  wire                                        mgr62__std__lane0_strm1_data_valid  ,

            // manager 62, lane 1, stream 0      
            input   wire                                        std__mgr62__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane1_strm0_data        ,
            output  wire                                        mgr62__std__lane1_strm0_data_valid  ,

            // manager 62, lane 1, stream 1      
            input   wire                                        std__mgr62__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane1_strm1_data        ,
            output  wire                                        mgr62__std__lane1_strm1_data_valid  ,

            // manager 62, lane 2, stream 0      
            input   wire                                        std__mgr62__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane2_strm0_data        ,
            output  wire                                        mgr62__std__lane2_strm0_data_valid  ,

            // manager 62, lane 2, stream 1      
            input   wire                                        std__mgr62__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane2_strm1_data        ,
            output  wire                                        mgr62__std__lane2_strm1_data_valid  ,

            // manager 62, lane 3, stream 0      
            input   wire                                        std__mgr62__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane3_strm0_data        ,
            output  wire                                        mgr62__std__lane3_strm0_data_valid  ,

            // manager 62, lane 3, stream 1      
            input   wire                                        std__mgr62__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane3_strm1_data        ,
            output  wire                                        mgr62__std__lane3_strm1_data_valid  ,

            // manager 62, lane 4, stream 0      
            input   wire                                        std__mgr62__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane4_strm0_data        ,
            output  wire                                        mgr62__std__lane4_strm0_data_valid  ,

            // manager 62, lane 4, stream 1      
            input   wire                                        std__mgr62__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane4_strm1_data        ,
            output  wire                                        mgr62__std__lane4_strm1_data_valid  ,

            // manager 62, lane 5, stream 0      
            input   wire                                        std__mgr62__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane5_strm0_data        ,
            output  wire                                        mgr62__std__lane5_strm0_data_valid  ,

            // manager 62, lane 5, stream 1      
            input   wire                                        std__mgr62__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane5_strm1_data        ,
            output  wire                                        mgr62__std__lane5_strm1_data_valid  ,

            // manager 62, lane 6, stream 0      
            input   wire                                        std__mgr62__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane6_strm0_data        ,
            output  wire                                        mgr62__std__lane6_strm0_data_valid  ,

            // manager 62, lane 6, stream 1      
            input   wire                                        std__mgr62__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane6_strm1_data        ,
            output  wire                                        mgr62__std__lane6_strm1_data_valid  ,

            // manager 62, lane 7, stream 0      
            input   wire                                        std__mgr62__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane7_strm0_data        ,
            output  wire                                        mgr62__std__lane7_strm0_data_valid  ,

            // manager 62, lane 7, stream 1      
            input   wire                                        std__mgr62__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane7_strm1_data        ,
            output  wire                                        mgr62__std__lane7_strm1_data_valid  ,

            // manager 62, lane 8, stream 0      
            input   wire                                        std__mgr62__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane8_strm0_data        ,
            output  wire                                        mgr62__std__lane8_strm0_data_valid  ,

            // manager 62, lane 8, stream 1      
            input   wire                                        std__mgr62__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane8_strm1_data        ,
            output  wire                                        mgr62__std__lane8_strm1_data_valid  ,

            // manager 62, lane 9, stream 0      
            input   wire                                        std__mgr62__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane9_strm0_data        ,
            output  wire                                        mgr62__std__lane9_strm0_data_valid  ,

            // manager 62, lane 9, stream 1      
            input   wire                                        std__mgr62__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane9_strm1_data        ,
            output  wire                                        mgr62__std__lane9_strm1_data_valid  ,

            // manager 62, lane 10, stream 0      
            input   wire                                        std__mgr62__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane10_strm0_data        ,
            output  wire                                        mgr62__std__lane10_strm0_data_valid  ,

            // manager 62, lane 10, stream 1      
            input   wire                                        std__mgr62__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane10_strm1_data        ,
            output  wire                                        mgr62__std__lane10_strm1_data_valid  ,

            // manager 62, lane 11, stream 0      
            input   wire                                        std__mgr62__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane11_strm0_data        ,
            output  wire                                        mgr62__std__lane11_strm0_data_valid  ,

            // manager 62, lane 11, stream 1      
            input   wire                                        std__mgr62__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane11_strm1_data        ,
            output  wire                                        mgr62__std__lane11_strm1_data_valid  ,

            // manager 62, lane 12, stream 0      
            input   wire                                        std__mgr62__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane12_strm0_data        ,
            output  wire                                        mgr62__std__lane12_strm0_data_valid  ,

            // manager 62, lane 12, stream 1      
            input   wire                                        std__mgr62__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane12_strm1_data        ,
            output  wire                                        mgr62__std__lane12_strm1_data_valid  ,

            // manager 62, lane 13, stream 0      
            input   wire                                        std__mgr62__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane13_strm0_data        ,
            output  wire                                        mgr62__std__lane13_strm0_data_valid  ,

            // manager 62, lane 13, stream 1      
            input   wire                                        std__mgr62__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane13_strm1_data        ,
            output  wire                                        mgr62__std__lane13_strm1_data_valid  ,

            // manager 62, lane 14, stream 0      
            input   wire                                        std__mgr62__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane14_strm0_data        ,
            output  wire                                        mgr62__std__lane14_strm0_data_valid  ,

            // manager 62, lane 14, stream 1      
            input   wire                                        std__mgr62__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane14_strm1_data        ,
            output  wire                                        mgr62__std__lane14_strm1_data_valid  ,

            // manager 62, lane 15, stream 0      
            input   wire                                        std__mgr62__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane15_strm0_data        ,
            output  wire                                        mgr62__std__lane15_strm0_data_valid  ,

            // manager 62, lane 15, stream 1      
            input   wire                                        std__mgr62__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane15_strm1_data        ,
            output  wire                                        mgr62__std__lane15_strm1_data_valid  ,

            // manager 62, lane 16, stream 0      
            input   wire                                        std__mgr62__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane16_strm0_data        ,
            output  wire                                        mgr62__std__lane16_strm0_data_valid  ,

            // manager 62, lane 16, stream 1      
            input   wire                                        std__mgr62__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane16_strm1_data        ,
            output  wire                                        mgr62__std__lane16_strm1_data_valid  ,

            // manager 62, lane 17, stream 0      
            input   wire                                        std__mgr62__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane17_strm0_data        ,
            output  wire                                        mgr62__std__lane17_strm0_data_valid  ,

            // manager 62, lane 17, stream 1      
            input   wire                                        std__mgr62__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane17_strm1_data        ,
            output  wire                                        mgr62__std__lane17_strm1_data_valid  ,

            // manager 62, lane 18, stream 0      
            input   wire                                        std__mgr62__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane18_strm0_data        ,
            output  wire                                        mgr62__std__lane18_strm0_data_valid  ,

            // manager 62, lane 18, stream 1      
            input   wire                                        std__mgr62__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane18_strm1_data        ,
            output  wire                                        mgr62__std__lane18_strm1_data_valid  ,

            // manager 62, lane 19, stream 0      
            input   wire                                        std__mgr62__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane19_strm0_data        ,
            output  wire                                        mgr62__std__lane19_strm0_data_valid  ,

            // manager 62, lane 19, stream 1      
            input   wire                                        std__mgr62__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane19_strm1_data        ,
            output  wire                                        mgr62__std__lane19_strm1_data_valid  ,

            // manager 62, lane 20, stream 0      
            input   wire                                        std__mgr62__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane20_strm0_data        ,
            output  wire                                        mgr62__std__lane20_strm0_data_valid  ,

            // manager 62, lane 20, stream 1      
            input   wire                                        std__mgr62__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane20_strm1_data        ,
            output  wire                                        mgr62__std__lane20_strm1_data_valid  ,

            // manager 62, lane 21, stream 0      
            input   wire                                        std__mgr62__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane21_strm0_data        ,
            output  wire                                        mgr62__std__lane21_strm0_data_valid  ,

            // manager 62, lane 21, stream 1      
            input   wire                                        std__mgr62__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane21_strm1_data        ,
            output  wire                                        mgr62__std__lane21_strm1_data_valid  ,

            // manager 62, lane 22, stream 0      
            input   wire                                        std__mgr62__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane22_strm0_data        ,
            output  wire                                        mgr62__std__lane22_strm0_data_valid  ,

            // manager 62, lane 22, stream 1      
            input   wire                                        std__mgr62__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane22_strm1_data        ,
            output  wire                                        mgr62__std__lane22_strm1_data_valid  ,

            // manager 62, lane 23, stream 0      
            input   wire                                        std__mgr62__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane23_strm0_data        ,
            output  wire                                        mgr62__std__lane23_strm0_data_valid  ,

            // manager 62, lane 23, stream 1      
            input   wire                                        std__mgr62__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane23_strm1_data        ,
            output  wire                                        mgr62__std__lane23_strm1_data_valid  ,

            // manager 62, lane 24, stream 0      
            input   wire                                        std__mgr62__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane24_strm0_data        ,
            output  wire                                        mgr62__std__lane24_strm0_data_valid  ,

            // manager 62, lane 24, stream 1      
            input   wire                                        std__mgr62__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane24_strm1_data        ,
            output  wire                                        mgr62__std__lane24_strm1_data_valid  ,

            // manager 62, lane 25, stream 0      
            input   wire                                        std__mgr62__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane25_strm0_data        ,
            output  wire                                        mgr62__std__lane25_strm0_data_valid  ,

            // manager 62, lane 25, stream 1      
            input   wire                                        std__mgr62__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane25_strm1_data        ,
            output  wire                                        mgr62__std__lane25_strm1_data_valid  ,

            // manager 62, lane 26, stream 0      
            input   wire                                        std__mgr62__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane26_strm0_data        ,
            output  wire                                        mgr62__std__lane26_strm0_data_valid  ,

            // manager 62, lane 26, stream 1      
            input   wire                                        std__mgr62__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane26_strm1_data        ,
            output  wire                                        mgr62__std__lane26_strm1_data_valid  ,

            // manager 62, lane 27, stream 0      
            input   wire                                        std__mgr62__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane27_strm0_data        ,
            output  wire                                        mgr62__std__lane27_strm0_data_valid  ,

            // manager 62, lane 27, stream 1      
            input   wire                                        std__mgr62__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane27_strm1_data        ,
            output  wire                                        mgr62__std__lane27_strm1_data_valid  ,

            // manager 62, lane 28, stream 0      
            input   wire                                        std__mgr62__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane28_strm0_data        ,
            output  wire                                        mgr62__std__lane28_strm0_data_valid  ,

            // manager 62, lane 28, stream 1      
            input   wire                                        std__mgr62__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane28_strm1_data        ,
            output  wire                                        mgr62__std__lane28_strm1_data_valid  ,

            // manager 62, lane 29, stream 0      
            input   wire                                        std__mgr62__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane29_strm0_data        ,
            output  wire                                        mgr62__std__lane29_strm0_data_valid  ,

            // manager 62, lane 29, stream 1      
            input   wire                                        std__mgr62__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane29_strm1_data        ,
            output  wire                                        mgr62__std__lane29_strm1_data_valid  ,

            // manager 62, lane 30, stream 0      
            input   wire                                        std__mgr62__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane30_strm0_data        ,
            output  wire                                        mgr62__std__lane30_strm0_data_valid  ,

            // manager 62, lane 30, stream 1      
            input   wire                                        std__mgr62__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane30_strm1_data        ,
            output  wire                                        mgr62__std__lane30_strm1_data_valid  ,

            // manager 62, lane 31, stream 0      
            input   wire                                        std__mgr62__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane31_strm0_data        ,
            output  wire                                        mgr62__std__lane31_strm0_data_valid  ,

            // manager 62, lane 31, stream 1      
            input   wire                                        std__mgr62__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr62__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr62__std__lane31_strm1_data        ,
            output  wire                                        mgr62__std__lane31_strm1_data_valid  ,

            //-----------------------------------------------------------
            // Manager Lane arguments to the PE                          

            // manager 63, lane 0, stream 0      
            input   wire                                        std__mgr63__lane0_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane0_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane0_strm0_data        ,
            output  wire                                        mgr63__std__lane0_strm0_data_valid  ,

            // manager 63, lane 0, stream 1      
            input   wire                                        std__mgr63__lane0_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane0_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane0_strm1_data        ,
            output  wire                                        mgr63__std__lane0_strm1_data_valid  ,

            // manager 63, lane 1, stream 0      
            input   wire                                        std__mgr63__lane1_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane1_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane1_strm0_data        ,
            output  wire                                        mgr63__std__lane1_strm0_data_valid  ,

            // manager 63, lane 1, stream 1      
            input   wire                                        std__mgr63__lane1_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane1_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane1_strm1_data        ,
            output  wire                                        mgr63__std__lane1_strm1_data_valid  ,

            // manager 63, lane 2, stream 0      
            input   wire                                        std__mgr63__lane2_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane2_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane2_strm0_data        ,
            output  wire                                        mgr63__std__lane2_strm0_data_valid  ,

            // manager 63, lane 2, stream 1      
            input   wire                                        std__mgr63__lane2_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane2_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane2_strm1_data        ,
            output  wire                                        mgr63__std__lane2_strm1_data_valid  ,

            // manager 63, lane 3, stream 0      
            input   wire                                        std__mgr63__lane3_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane3_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane3_strm0_data        ,
            output  wire                                        mgr63__std__lane3_strm0_data_valid  ,

            // manager 63, lane 3, stream 1      
            input   wire                                        std__mgr63__lane3_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane3_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane3_strm1_data        ,
            output  wire                                        mgr63__std__lane3_strm1_data_valid  ,

            // manager 63, lane 4, stream 0      
            input   wire                                        std__mgr63__lane4_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane4_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane4_strm0_data        ,
            output  wire                                        mgr63__std__lane4_strm0_data_valid  ,

            // manager 63, lane 4, stream 1      
            input   wire                                        std__mgr63__lane4_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane4_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane4_strm1_data        ,
            output  wire                                        mgr63__std__lane4_strm1_data_valid  ,

            // manager 63, lane 5, stream 0      
            input   wire                                        std__mgr63__lane5_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane5_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane5_strm0_data        ,
            output  wire                                        mgr63__std__lane5_strm0_data_valid  ,

            // manager 63, lane 5, stream 1      
            input   wire                                        std__mgr63__lane5_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane5_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane5_strm1_data        ,
            output  wire                                        mgr63__std__lane5_strm1_data_valid  ,

            // manager 63, lane 6, stream 0      
            input   wire                                        std__mgr63__lane6_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane6_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane6_strm0_data        ,
            output  wire                                        mgr63__std__lane6_strm0_data_valid  ,

            // manager 63, lane 6, stream 1      
            input   wire                                        std__mgr63__lane6_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane6_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane6_strm1_data        ,
            output  wire                                        mgr63__std__lane6_strm1_data_valid  ,

            // manager 63, lane 7, stream 0      
            input   wire                                        std__mgr63__lane7_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane7_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane7_strm0_data        ,
            output  wire                                        mgr63__std__lane7_strm0_data_valid  ,

            // manager 63, lane 7, stream 1      
            input   wire                                        std__mgr63__lane7_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane7_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane7_strm1_data        ,
            output  wire                                        mgr63__std__lane7_strm1_data_valid  ,

            // manager 63, lane 8, stream 0      
            input   wire                                        std__mgr63__lane8_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane8_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane8_strm0_data        ,
            output  wire                                        mgr63__std__lane8_strm0_data_valid  ,

            // manager 63, lane 8, stream 1      
            input   wire                                        std__mgr63__lane8_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane8_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane8_strm1_data        ,
            output  wire                                        mgr63__std__lane8_strm1_data_valid  ,

            // manager 63, lane 9, stream 0      
            input   wire                                        std__mgr63__lane9_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane9_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane9_strm0_data        ,
            output  wire                                        mgr63__std__lane9_strm0_data_valid  ,

            // manager 63, lane 9, stream 1      
            input   wire                                        std__mgr63__lane9_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane9_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane9_strm1_data        ,
            output  wire                                        mgr63__std__lane9_strm1_data_valid  ,

            // manager 63, lane 10, stream 0      
            input   wire                                        std__mgr63__lane10_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane10_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane10_strm0_data        ,
            output  wire                                        mgr63__std__lane10_strm0_data_valid  ,

            // manager 63, lane 10, stream 1      
            input   wire                                        std__mgr63__lane10_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane10_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane10_strm1_data        ,
            output  wire                                        mgr63__std__lane10_strm1_data_valid  ,

            // manager 63, lane 11, stream 0      
            input   wire                                        std__mgr63__lane11_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane11_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane11_strm0_data        ,
            output  wire                                        mgr63__std__lane11_strm0_data_valid  ,

            // manager 63, lane 11, stream 1      
            input   wire                                        std__mgr63__lane11_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane11_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane11_strm1_data        ,
            output  wire                                        mgr63__std__lane11_strm1_data_valid  ,

            // manager 63, lane 12, stream 0      
            input   wire                                        std__mgr63__lane12_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane12_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane12_strm0_data        ,
            output  wire                                        mgr63__std__lane12_strm0_data_valid  ,

            // manager 63, lane 12, stream 1      
            input   wire                                        std__mgr63__lane12_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane12_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane12_strm1_data        ,
            output  wire                                        mgr63__std__lane12_strm1_data_valid  ,

            // manager 63, lane 13, stream 0      
            input   wire                                        std__mgr63__lane13_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane13_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane13_strm0_data        ,
            output  wire                                        mgr63__std__lane13_strm0_data_valid  ,

            // manager 63, lane 13, stream 1      
            input   wire                                        std__mgr63__lane13_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane13_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane13_strm1_data        ,
            output  wire                                        mgr63__std__lane13_strm1_data_valid  ,

            // manager 63, lane 14, stream 0      
            input   wire                                        std__mgr63__lane14_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane14_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane14_strm0_data        ,
            output  wire                                        mgr63__std__lane14_strm0_data_valid  ,

            // manager 63, lane 14, stream 1      
            input   wire                                        std__mgr63__lane14_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane14_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane14_strm1_data        ,
            output  wire                                        mgr63__std__lane14_strm1_data_valid  ,

            // manager 63, lane 15, stream 0      
            input   wire                                        std__mgr63__lane15_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane15_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane15_strm0_data        ,
            output  wire                                        mgr63__std__lane15_strm0_data_valid  ,

            // manager 63, lane 15, stream 1      
            input   wire                                        std__mgr63__lane15_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane15_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane15_strm1_data        ,
            output  wire                                        mgr63__std__lane15_strm1_data_valid  ,

            // manager 63, lane 16, stream 0      
            input   wire                                        std__mgr63__lane16_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane16_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane16_strm0_data        ,
            output  wire                                        mgr63__std__lane16_strm0_data_valid  ,

            // manager 63, lane 16, stream 1      
            input   wire                                        std__mgr63__lane16_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane16_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane16_strm1_data        ,
            output  wire                                        mgr63__std__lane16_strm1_data_valid  ,

            // manager 63, lane 17, stream 0      
            input   wire                                        std__mgr63__lane17_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane17_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane17_strm0_data        ,
            output  wire                                        mgr63__std__lane17_strm0_data_valid  ,

            // manager 63, lane 17, stream 1      
            input   wire                                        std__mgr63__lane17_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane17_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane17_strm1_data        ,
            output  wire                                        mgr63__std__lane17_strm1_data_valid  ,

            // manager 63, lane 18, stream 0      
            input   wire                                        std__mgr63__lane18_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane18_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane18_strm0_data        ,
            output  wire                                        mgr63__std__lane18_strm0_data_valid  ,

            // manager 63, lane 18, stream 1      
            input   wire                                        std__mgr63__lane18_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane18_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane18_strm1_data        ,
            output  wire                                        mgr63__std__lane18_strm1_data_valid  ,

            // manager 63, lane 19, stream 0      
            input   wire                                        std__mgr63__lane19_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane19_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane19_strm0_data        ,
            output  wire                                        mgr63__std__lane19_strm0_data_valid  ,

            // manager 63, lane 19, stream 1      
            input   wire                                        std__mgr63__lane19_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane19_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane19_strm1_data        ,
            output  wire                                        mgr63__std__lane19_strm1_data_valid  ,

            // manager 63, lane 20, stream 0      
            input   wire                                        std__mgr63__lane20_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane20_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane20_strm0_data        ,
            output  wire                                        mgr63__std__lane20_strm0_data_valid  ,

            // manager 63, lane 20, stream 1      
            input   wire                                        std__mgr63__lane20_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane20_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane20_strm1_data        ,
            output  wire                                        mgr63__std__lane20_strm1_data_valid  ,

            // manager 63, lane 21, stream 0      
            input   wire                                        std__mgr63__lane21_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane21_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane21_strm0_data        ,
            output  wire                                        mgr63__std__lane21_strm0_data_valid  ,

            // manager 63, lane 21, stream 1      
            input   wire                                        std__mgr63__lane21_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane21_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane21_strm1_data        ,
            output  wire                                        mgr63__std__lane21_strm1_data_valid  ,

            // manager 63, lane 22, stream 0      
            input   wire                                        std__mgr63__lane22_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane22_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane22_strm0_data        ,
            output  wire                                        mgr63__std__lane22_strm0_data_valid  ,

            // manager 63, lane 22, stream 1      
            input   wire                                        std__mgr63__lane22_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane22_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane22_strm1_data        ,
            output  wire                                        mgr63__std__lane22_strm1_data_valid  ,

            // manager 63, lane 23, stream 0      
            input   wire                                        std__mgr63__lane23_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane23_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane23_strm0_data        ,
            output  wire                                        mgr63__std__lane23_strm0_data_valid  ,

            // manager 63, lane 23, stream 1      
            input   wire                                        std__mgr63__lane23_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane23_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane23_strm1_data        ,
            output  wire                                        mgr63__std__lane23_strm1_data_valid  ,

            // manager 63, lane 24, stream 0      
            input   wire                                        std__mgr63__lane24_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane24_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane24_strm0_data        ,
            output  wire                                        mgr63__std__lane24_strm0_data_valid  ,

            // manager 63, lane 24, stream 1      
            input   wire                                        std__mgr63__lane24_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane24_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane24_strm1_data        ,
            output  wire                                        mgr63__std__lane24_strm1_data_valid  ,

            // manager 63, lane 25, stream 0      
            input   wire                                        std__mgr63__lane25_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane25_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane25_strm0_data        ,
            output  wire                                        mgr63__std__lane25_strm0_data_valid  ,

            // manager 63, lane 25, stream 1      
            input   wire                                        std__mgr63__lane25_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane25_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane25_strm1_data        ,
            output  wire                                        mgr63__std__lane25_strm1_data_valid  ,

            // manager 63, lane 26, stream 0      
            input   wire                                        std__mgr63__lane26_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane26_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane26_strm0_data        ,
            output  wire                                        mgr63__std__lane26_strm0_data_valid  ,

            // manager 63, lane 26, stream 1      
            input   wire                                        std__mgr63__lane26_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane26_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane26_strm1_data        ,
            output  wire                                        mgr63__std__lane26_strm1_data_valid  ,

            // manager 63, lane 27, stream 0      
            input   wire                                        std__mgr63__lane27_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane27_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane27_strm0_data        ,
            output  wire                                        mgr63__std__lane27_strm0_data_valid  ,

            // manager 63, lane 27, stream 1      
            input   wire                                        std__mgr63__lane27_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane27_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane27_strm1_data        ,
            output  wire                                        mgr63__std__lane27_strm1_data_valid  ,

            // manager 63, lane 28, stream 0      
            input   wire                                        std__mgr63__lane28_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane28_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane28_strm0_data        ,
            output  wire                                        mgr63__std__lane28_strm0_data_valid  ,

            // manager 63, lane 28, stream 1      
            input   wire                                        std__mgr63__lane28_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane28_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane28_strm1_data        ,
            output  wire                                        mgr63__std__lane28_strm1_data_valid  ,

            // manager 63, lane 29, stream 0      
            input   wire                                        std__mgr63__lane29_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane29_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane29_strm0_data        ,
            output  wire                                        mgr63__std__lane29_strm0_data_valid  ,

            // manager 63, lane 29, stream 1      
            input   wire                                        std__mgr63__lane29_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane29_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane29_strm1_data        ,
            output  wire                                        mgr63__std__lane29_strm1_data_valid  ,

            // manager 63, lane 30, stream 0      
            input   wire                                        std__mgr63__lane30_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane30_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane30_strm0_data        ,
            output  wire                                        mgr63__std__lane30_strm0_data_valid  ,

            // manager 63, lane 30, stream 1      
            input   wire                                        std__mgr63__lane30_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane30_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane30_strm1_data        ,
            output  wire                                        mgr63__std__lane30_strm1_data_valid  ,

            // manager 63, lane 31, stream 0      
            input   wire                                        std__mgr63__lane31_strm0_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane31_strm0_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane31_strm0_data        ,
            output  wire                                        mgr63__std__lane31_strm0_data_valid  ,

            // manager 63, lane 31, stream 1      
            input   wire                                        std__mgr63__lane31_strm1_ready       ,
            output  wire  [`COMMON_STD_INTF_CNTL_RANGE      ]   mgr63__std__lane31_strm1_cntl        ,
            output  wire  [`STACK_DOWN_INTF_STRM_DATA_RANGE ]   mgr63__std__lane31_strm1_data        ,
            output  wire                                        mgr63__std__lane31_strm1_data_valid  ,
