
            begin
              wait(final_operation[0].triggered) ; // we start waiting before the event will occur
              //@(final_operation[0]) ;
              //$display("@%0t LEE: Received final operation event for manager 0\n", $time);
            end
            begin
              wait(final_operation[1].triggered) ; // we start waiting before the event will occur
              //@(final_operation[1]) ;
              //$display("@%0t LEE: Received final operation event for manager 1\n", $time);
            end
            begin
              wait(final_operation[2].triggered) ; // we start waiting before the event will occur
              //@(final_operation[2]) ;
              //$display("@%0t LEE: Received final operation event for manager 2\n", $time);
            end
            begin
              wait(final_operation[3].triggered) ; // we start waiting before the event will occur
              //@(final_operation[3]) ;
              //$display("@%0t LEE: Received final operation event for manager 3\n", $time);
            end
            begin
              wait(final_operation[4].triggered) ; // we start waiting before the event will occur
              //@(final_operation[4]) ;
              //$display("@%0t LEE: Received final operation event for manager 4\n", $time);
            end
            begin
              wait(final_operation[5].triggered) ; // we start waiting before the event will occur
              //@(final_operation[5]) ;
              //$display("@%0t LEE: Received final operation event for manager 5\n", $time);
            end
            begin
              wait(final_operation[6].triggered) ; // we start waiting before the event will occur
              //@(final_operation[6]) ;
              //$display("@%0t LEE: Received final operation event for manager 6\n", $time);
            end
            begin
              wait(final_operation[7].triggered) ; // we start waiting before the event will occur
              //@(final_operation[7]) ;
              //$display("@%0t LEE: Received final operation event for manager 7\n", $time);
            end
            begin
              wait(final_operation[8].triggered) ; // we start waiting before the event will occur
              //@(final_operation[8]) ;
              //$display("@%0t LEE: Received final operation event for manager 8\n", $time);
            end
            begin
              wait(final_operation[9].triggered) ; // we start waiting before the event will occur
              //@(final_operation[9]) ;
              //$display("@%0t LEE: Received final operation event for manager 9\n", $time);
            end
            begin
              wait(final_operation[10].triggered) ; // we start waiting before the event will occur
              //@(final_operation[10]) ;
              //$display("@%0t LEE: Received final operation event for manager 10\n", $time);
            end
            begin
              wait(final_operation[11].triggered) ; // we start waiting before the event will occur
              //@(final_operation[11]) ;
              //$display("@%0t LEE: Received final operation event for manager 11\n", $time);
            end
            begin
              wait(final_operation[12].triggered) ; // we start waiting before the event will occur
              //@(final_operation[12]) ;
              //$display("@%0t LEE: Received final operation event for manager 12\n", $time);
            end
            begin
              wait(final_operation[13].triggered) ; // we start waiting before the event will occur
              //@(final_operation[13]) ;
              //$display("@%0t LEE: Received final operation event for manager 13\n", $time);
            end
            begin
              wait(final_operation[14].triggered) ; // we start waiting before the event will occur
              //@(final_operation[14]) ;
              //$display("@%0t LEE: Received final operation event for manager 14\n", $time);
            end
            begin
              wait(final_operation[15].triggered) ; // we start waiting before the event will occur
              //@(final_operation[15]) ;
              //$display("@%0t LEE: Received final operation event for manager 15\n", $time);
            end
            begin
              wait(final_operation[16].triggered) ; // we start waiting before the event will occur
              //@(final_operation[16]) ;
              //$display("@%0t LEE: Received final operation event for manager 16\n", $time);
            end
            begin
              wait(final_operation[17].triggered) ; // we start waiting before the event will occur
              //@(final_operation[17]) ;
              //$display("@%0t LEE: Received final operation event for manager 17\n", $time);
            end
            begin
              wait(final_operation[18].triggered) ; // we start waiting before the event will occur
              //@(final_operation[18]) ;
              //$display("@%0t LEE: Received final operation event for manager 18\n", $time);
            end
            begin
              wait(final_operation[19].triggered) ; // we start waiting before the event will occur
              //@(final_operation[19]) ;
              //$display("@%0t LEE: Received final operation event for manager 19\n", $time);
            end
            begin
              wait(final_operation[20].triggered) ; // we start waiting before the event will occur
              //@(final_operation[20]) ;
              //$display("@%0t LEE: Received final operation event for manager 20\n", $time);
            end
            begin
              wait(final_operation[21].triggered) ; // we start waiting before the event will occur
              //@(final_operation[21]) ;
              //$display("@%0t LEE: Received final operation event for manager 21\n", $time);
            end
            begin
              wait(final_operation[22].triggered) ; // we start waiting before the event will occur
              //@(final_operation[22]) ;
              //$display("@%0t LEE: Received final operation event for manager 22\n", $time);
            end
            begin
              wait(final_operation[23].triggered) ; // we start waiting before the event will occur
              //@(final_operation[23]) ;
              //$display("@%0t LEE: Received final operation event for manager 23\n", $time);
            end
            begin
              wait(final_operation[24].triggered) ; // we start waiting before the event will occur
              //@(final_operation[24]) ;
              //$display("@%0t LEE: Received final operation event for manager 24\n", $time);
            end
            begin
              wait(final_operation[25].triggered) ; // we start waiting before the event will occur
              //@(final_operation[25]) ;
              //$display("@%0t LEE: Received final operation event for manager 25\n", $time);
            end
            begin
              wait(final_operation[26].triggered) ; // we start waiting before the event will occur
              //@(final_operation[26]) ;
              //$display("@%0t LEE: Received final operation event for manager 26\n", $time);
            end
            begin
              wait(final_operation[27].triggered) ; // we start waiting before the event will occur
              //@(final_operation[27]) ;
              //$display("@%0t LEE: Received final operation event for manager 27\n", $time);
            end
            begin
              wait(final_operation[28].triggered) ; // we start waiting before the event will occur
              //@(final_operation[28]) ;
              //$display("@%0t LEE: Received final operation event for manager 28\n", $time);
            end
            begin
              wait(final_operation[29].triggered) ; // we start waiting before the event will occur
              //@(final_operation[29]) ;
              //$display("@%0t LEE: Received final operation event for manager 29\n", $time);
            end
            begin
              wait(final_operation[30].triggered) ; // we start waiting before the event will occur
              //@(final_operation[30]) ;
              //$display("@%0t LEE: Received final operation event for manager 30\n", $time);
            end
            begin
              wait(final_operation[31].triggered) ; // we start waiting before the event will occur
              //@(final_operation[31]) ;
              //$display("@%0t LEE: Received final operation event for manager 31\n", $time);
            end
            begin
              wait(final_operation[32].triggered) ; // we start waiting before the event will occur
              //@(final_operation[32]) ;
              //$display("@%0t LEE: Received final operation event for manager 32\n", $time);
            end
            begin
              wait(final_operation[33].triggered) ; // we start waiting before the event will occur
              //@(final_operation[33]) ;
              //$display("@%0t LEE: Received final operation event for manager 33\n", $time);
            end
            begin
              wait(final_operation[34].triggered) ; // we start waiting before the event will occur
              //@(final_operation[34]) ;
              //$display("@%0t LEE: Received final operation event for manager 34\n", $time);
            end
            begin
              wait(final_operation[35].triggered) ; // we start waiting before the event will occur
              //@(final_operation[35]) ;
              //$display("@%0t LEE: Received final operation event for manager 35\n", $time);
            end
            begin
              wait(final_operation[36].triggered) ; // we start waiting before the event will occur
              //@(final_operation[36]) ;
              //$display("@%0t LEE: Received final operation event for manager 36\n", $time);
            end
            begin
              wait(final_operation[37].triggered) ; // we start waiting before the event will occur
              //@(final_operation[37]) ;
              //$display("@%0t LEE: Received final operation event for manager 37\n", $time);
            end
            begin
              wait(final_operation[38].triggered) ; // we start waiting before the event will occur
              //@(final_operation[38]) ;
              //$display("@%0t LEE: Received final operation event for manager 38\n", $time);
            end
            begin
              wait(final_operation[39].triggered) ; // we start waiting before the event will occur
              //@(final_operation[39]) ;
              //$display("@%0t LEE: Received final operation event for manager 39\n", $time);
            end
            begin
              wait(final_operation[40].triggered) ; // we start waiting before the event will occur
              //@(final_operation[40]) ;
              //$display("@%0t LEE: Received final operation event for manager 40\n", $time);
            end
            begin
              wait(final_operation[41].triggered) ; // we start waiting before the event will occur
              //@(final_operation[41]) ;
              //$display("@%0t LEE: Received final operation event for manager 41\n", $time);
            end
            begin
              wait(final_operation[42].triggered) ; // we start waiting before the event will occur
              //@(final_operation[42]) ;
              //$display("@%0t LEE: Received final operation event for manager 42\n", $time);
            end
            begin
              wait(final_operation[43].triggered) ; // we start waiting before the event will occur
              //@(final_operation[43]) ;
              //$display("@%0t LEE: Received final operation event for manager 43\n", $time);
            end
            begin
              wait(final_operation[44].triggered) ; // we start waiting before the event will occur
              //@(final_operation[44]) ;
              //$display("@%0t LEE: Received final operation event for manager 44\n", $time);
            end
            begin
              wait(final_operation[45].triggered) ; // we start waiting before the event will occur
              //@(final_operation[45]) ;
              //$display("@%0t LEE: Received final operation event for manager 45\n", $time);
            end
            begin
              wait(final_operation[46].triggered) ; // we start waiting before the event will occur
              //@(final_operation[46]) ;
              //$display("@%0t LEE: Received final operation event for manager 46\n", $time);
            end
            begin
              wait(final_operation[47].triggered) ; // we start waiting before the event will occur
              //@(final_operation[47]) ;
              //$display("@%0t LEE: Received final operation event for manager 47\n", $time);
            end
            begin
              wait(final_operation[48].triggered) ; // we start waiting before the event will occur
              //@(final_operation[48]) ;
              //$display("@%0t LEE: Received final operation event for manager 48\n", $time);
            end
            begin
              wait(final_operation[49].triggered) ; // we start waiting before the event will occur
              //@(final_operation[49]) ;
              //$display("@%0t LEE: Received final operation event for manager 49\n", $time);
            end
            begin
              wait(final_operation[50].triggered) ; // we start waiting before the event will occur
              //@(final_operation[50]) ;
              //$display("@%0t LEE: Received final operation event for manager 50\n", $time);
            end
            begin
              wait(final_operation[51].triggered) ; // we start waiting before the event will occur
              //@(final_operation[51]) ;
              //$display("@%0t LEE: Received final operation event for manager 51\n", $time);
            end
            begin
              wait(final_operation[52].triggered) ; // we start waiting before the event will occur
              //@(final_operation[52]) ;
              //$display("@%0t LEE: Received final operation event for manager 52\n", $time);
            end
            begin
              wait(final_operation[53].triggered) ; // we start waiting before the event will occur
              //@(final_operation[53]) ;
              //$display("@%0t LEE: Received final operation event for manager 53\n", $time);
            end
            begin
              wait(final_operation[54].triggered) ; // we start waiting before the event will occur
              //@(final_operation[54]) ;
              //$display("@%0t LEE: Received final operation event for manager 54\n", $time);
            end
            begin
              wait(final_operation[55].triggered) ; // we start waiting before the event will occur
              //@(final_operation[55]) ;
              //$display("@%0t LEE: Received final operation event for manager 55\n", $time);
            end
            begin
              wait(final_operation[56].triggered) ; // we start waiting before the event will occur
              //@(final_operation[56]) ;
              //$display("@%0t LEE: Received final operation event for manager 56\n", $time);
            end
            begin
              wait(final_operation[57].triggered) ; // we start waiting before the event will occur
              //@(final_operation[57]) ;
              //$display("@%0t LEE: Received final operation event for manager 57\n", $time);
            end
            begin
              wait(final_operation[58].triggered) ; // we start waiting before the event will occur
              //@(final_operation[58]) ;
              //$display("@%0t LEE: Received final operation event for manager 58\n", $time);
            end
            begin
              wait(final_operation[59].triggered) ; // we start waiting before the event will occur
              //@(final_operation[59]) ;
              //$display("@%0t LEE: Received final operation event for manager 59\n", $time);
            end
            begin
              wait(final_operation[60].triggered) ; // we start waiting before the event will occur
              //@(final_operation[60]) ;
              //$display("@%0t LEE: Received final operation event for manager 60\n", $time);
            end
            begin
              wait(final_operation[61].triggered) ; // we start waiting before the event will occur
              //@(final_operation[61]) ;
              //$display("@%0t LEE: Received final operation event for manager 61\n", $time);
            end
            begin
              wait(final_operation[62].triggered) ; // we start waiting before the event will occur
              //@(final_operation[62]) ;
              //$display("@%0t LEE: Received final operation event for manager 62\n", $time);
            end
            begin
              wait(final_operation[63].triggered) ; // we start waiting before the event will occur
              //@(final_operation[63]) ;
              //$display("@%0t LEE: Received final operation event for manager 63\n", $time);
            end
