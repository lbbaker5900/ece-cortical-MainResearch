
            // Common (Scalar) Register(s)                
            .cntl__simd__rs0         ( cntl__simd__rs0        ),
            .cntl__simd__rs1         ( cntl__simd__rs1        ),

            // Lane 31             
            .cntl__simd__lane_r128   ( cntl__simd__lane_r128  ),
            .cntl__simd__lane_r129   ( cntl__simd__lane_r129  ),
            .cntl__simd__lane_r130   ( cntl__simd__lane_r130  ),
            .cntl__simd__lane_r131   ( cntl__simd__lane_r131  ),
            .cntl__simd__lane_r132   ( cntl__simd__lane_r132  ),
            .cntl__simd__lane_r133   ( cntl__simd__lane_r133  ),
            .cntl__simd__lane_r134   ( cntl__simd__lane_r134  ),
            .cntl__simd__lane_r135   ( cntl__simd__lane_r135  ),
