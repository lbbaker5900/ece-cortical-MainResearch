
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[0].numberOfLanes < 0)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[0].put(sys_operation_lane_gen[0]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[0];                                       
                //  end                                                        
            join_none                                                        
                                                                             
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[1].numberOfLanes < 1)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[1].put(sys_operation_lane_gen[1]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[1];                                       
                //  end                                                        
            join_none                                                        
                                                                             
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[2].numberOfLanes < 2)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[2].put(sys_operation_lane_gen[2]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[2];                                       
                //  end                                                        
            join_none                                                        
                                                                             
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[3].numberOfLanes < 3)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[3].put(sys_operation_lane_gen[3]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[3];                                       
                //  end                                                        
            join_none                                                        
                                                                             
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[4].numberOfLanes < 4)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[4].put(sys_operation_lane_gen[4]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[4];                                       
                //  end                                                        
            join_none                                                        
                                                                             
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[5].numberOfLanes < 5)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[5].put(sys_operation_lane_gen[5]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[5];                                       
                //  end                                                        
            join_none                                                        
                                                                             
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[6].numberOfLanes < 6)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[6].put(sys_operation_lane_gen[6]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[6];                                       
                //  end                                                        
            join_none                                                        
                                                                             
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[7].numberOfLanes < 7)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[7].put(sys_operation_lane_gen[7]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[7];                                       
                //  end                                                        
            join_none                                                        
                                                                             
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[8].numberOfLanes < 8)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[8].put(sys_operation_lane_gen[8]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[8];                                       
                //  end                                                        
            join_none                                                        
                                                                             
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[9].numberOfLanes < 9)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[9].put(sys_operation_lane_gen[9]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[9];                                       
                //  end                                                        
            join_none                                                        
                                                                             
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[10].numberOfLanes < 10)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[10].put(sys_operation_lane_gen[10]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[10];                                       
                //  end                                                        
            join_none                                                        
                                                                             
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[11].numberOfLanes < 11)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[11].put(sys_operation_lane_gen[11]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[11];                                       
                //  end                                                        
            join_none                                                        
                                                                             
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[12].numberOfLanes < 12)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[12].put(sys_operation_lane_gen[12]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[12];                                       
                //  end                                                        
            join_none                                                        
                                                                             
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[13].numberOfLanes < 13)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[13].put(sys_operation_lane_gen[13]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[13];                                       
                //  end                                                        
            join_none                                                        
                                                                             
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[14].numberOfLanes < 14)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[14].put(sys_operation_lane_gen[14]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[14];                                       
                //  end                                                        
            join_none                                                        
                                                                             
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[15].numberOfLanes < 15)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[15].put(sys_operation_lane_gen[15]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[15];                                       
                //  end                                                        
            join_none                                                        
                                                                             
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[16].numberOfLanes < 16)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[16].put(sys_operation_lane_gen[16]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[16];                                       
                //  end                                                        
            join_none                                                        
                                                                             
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[17].numberOfLanes < 17)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[17].put(sys_operation_lane_gen[17]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[17];                                       
                //  end                                                        
            join_none                                                        
                                                                             
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[18].numberOfLanes < 18)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[18].put(sys_operation_lane_gen[18]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[18];                                       
                //  end                                                        
            join_none                                                        
                                                                             
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[19].numberOfLanes < 19)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[19].put(sys_operation_lane_gen[19]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[19];                                       
                //  end                                                        
            join_none                                                        
                                                                             
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[20].numberOfLanes < 20)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[20].put(sys_operation_lane_gen[20]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[20];                                       
                //  end                                                        
            join_none                                                        
                                                                             
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[21].numberOfLanes < 21)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[21].put(sys_operation_lane_gen[21]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[21];                                       
                //  end                                                        
            join_none                                                        
                                                                             
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[22].numberOfLanes < 22)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[22].put(sys_operation_lane_gen[22]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[22];                                       
                //  end                                                        
            join_none                                                        
                                                                             
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[23].numberOfLanes < 23)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[23].put(sys_operation_lane_gen[23]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[23];                                       
                //  end                                                        
            join_none                                                        
                                                                             
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[24].numberOfLanes < 24)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[24].put(sys_operation_lane_gen[24]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[24];                                       
                //  end                                                        
            join_none                                                        
                                                                             
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[25].numberOfLanes < 25)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[25].put(sys_operation_lane_gen[25]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[25];                                       
                //  end                                                        
            join_none                                                        
                                                                             
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[26].numberOfLanes < 26)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[26].put(sys_operation_lane_gen[26]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[26];                                       
                //  end                                                        
            join_none                                                        
                                                                             
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[27].numberOfLanes < 27)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[27].put(sys_operation_lane_gen[27]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[27];                                       
                //  end                                                        
            join_none                                                        
                                                                             
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[28].numberOfLanes < 28)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[28].put(sys_operation_lane_gen[28]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[28];                                       
                //  end                                                        
            join_none                                                        
                                                                             
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[29].numberOfLanes < 29)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[29].put(sys_operation_lane_gen[29]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[29];                                       
                //  end                                                        
            join_none                                                        
                                                                             
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[30].numberOfLanes < 30)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[30].put(sys_operation_lane_gen[30]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[30];                                       
                //  end                                                        
            join_none                                                        
                                                                             
            fork                                                                                                                                  
                //if (sys_operation_lane_gen[31].numberOfLanes < 31)         
                //  begin
                    // Send to driver                                        
                    mgr2gen[31].put(sys_operation_lane_gen[31]) ;          
                    // now wait for generator                                
                    @mgr2gen_ack[31];                                       
                //  end                                                        
            join_none                                                        
                                                                             
