
  assign stOp_lane[0].scntl__dma__operation    = scntl__sdp__lane0_dma_operation ;
  assign stOp_lane[1].scntl__dma__operation    = scntl__sdp__lane1_dma_operation ;
  assign stOp_lane[2].scntl__dma__operation    = scntl__sdp__lane2_dma_operation ;
  assign stOp_lane[3].scntl__dma__operation    = scntl__sdp__lane3_dma_operation ;
  assign stOp_lane[4].scntl__dma__operation    = scntl__sdp__lane4_dma_operation ;
  assign stOp_lane[5].scntl__dma__operation    = scntl__sdp__lane5_dma_operation ;
  assign stOp_lane[6].scntl__dma__operation    = scntl__sdp__lane6_dma_operation ;
  assign stOp_lane[7].scntl__dma__operation    = scntl__sdp__lane7_dma_operation ;
  assign stOp_lane[8].scntl__dma__operation    = scntl__sdp__lane8_dma_operation ;
  assign stOp_lane[9].scntl__dma__operation    = scntl__sdp__lane9_dma_operation ;
  assign stOp_lane[10].scntl__dma__operation    = scntl__sdp__lane10_dma_operation ;
  assign stOp_lane[11].scntl__dma__operation    = scntl__sdp__lane11_dma_operation ;
  assign stOp_lane[12].scntl__dma__operation    = scntl__sdp__lane12_dma_operation ;
  assign stOp_lane[13].scntl__dma__operation    = scntl__sdp__lane13_dma_operation ;
  assign stOp_lane[14].scntl__dma__operation    = scntl__sdp__lane14_dma_operation ;
  assign stOp_lane[15].scntl__dma__operation    = scntl__sdp__lane15_dma_operation ;
  assign stOp_lane[16].scntl__dma__operation    = scntl__sdp__lane16_dma_operation ;
  assign stOp_lane[17].scntl__dma__operation    = scntl__sdp__lane17_dma_operation ;
  assign stOp_lane[18].scntl__dma__operation    = scntl__sdp__lane18_dma_operation ;
  assign stOp_lane[19].scntl__dma__operation    = scntl__sdp__lane19_dma_operation ;
  assign stOp_lane[20].scntl__dma__operation    = scntl__sdp__lane20_dma_operation ;
  assign stOp_lane[21].scntl__dma__operation    = scntl__sdp__lane21_dma_operation ;
  assign stOp_lane[22].scntl__dma__operation    = scntl__sdp__lane22_dma_operation ;
  assign stOp_lane[23].scntl__dma__operation    = scntl__sdp__lane23_dma_operation ;
  assign stOp_lane[24].scntl__dma__operation    = scntl__sdp__lane24_dma_operation ;
  assign stOp_lane[25].scntl__dma__operation    = scntl__sdp__lane25_dma_operation ;
  assign stOp_lane[26].scntl__dma__operation    = scntl__sdp__lane26_dma_operation ;
  assign stOp_lane[27].scntl__dma__operation    = scntl__sdp__lane27_dma_operation ;
  assign stOp_lane[28].scntl__dma__operation    = scntl__sdp__lane28_dma_operation ;
  assign stOp_lane[29].scntl__dma__operation    = scntl__sdp__lane29_dma_operation ;
  assign stOp_lane[30].scntl__dma__operation    = scntl__sdp__lane30_dma_operation ;
  assign stOp_lane[31].scntl__dma__operation    = scntl__sdp__lane31_dma_operation ;

  assign stOp_lane[0].scntl__dma__strm0_read_enable         = scntl__sdp__lane0_strm0_read_enable            ;
  assign stOp_lane[0].scntl__dma__strm0_write_enable        = scntl__sdp__lane0_strm0_write_enable           ;
  assign sdp__scntl__lane0_strm0_read_ready                 = stOp_lane[0].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane0_strm0_write_ready                = stOp_lane[0].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane0_strm0_read_complete              = stOp_lane[0].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane0_strm0_write_complete             = stOp_lane[0].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[0].scntl__dma__strm0_read_start_address  = scntl__sdp__lane0_strm0_read_start_address     ;
  assign stOp_lane[0].scntl__dma__strm0_write_start_address = scntl__sdp__lane0_strm0_write_start_address    ;
  assign stOp_lane[0].scntl__dma__type0                     = scntl__sdp__lane0_type0                        ;
  assign stOp_lane[0].scntl__dma__num_of_types0             = scntl__sdp__lane0_num_of_types0                ;
  assign stOp_lane[1].scntl__dma__strm0_read_enable         = scntl__sdp__lane1_strm0_read_enable            ;
  assign stOp_lane[1].scntl__dma__strm0_write_enable        = scntl__sdp__lane1_strm0_write_enable           ;
  assign sdp__scntl__lane1_strm0_read_ready                 = stOp_lane[1].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane1_strm0_write_ready                = stOp_lane[1].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane1_strm0_read_complete              = stOp_lane[1].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane1_strm0_write_complete             = stOp_lane[1].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[1].scntl__dma__strm0_read_start_address  = scntl__sdp__lane1_strm0_read_start_address     ;
  assign stOp_lane[1].scntl__dma__strm0_write_start_address = scntl__sdp__lane1_strm0_write_start_address    ;
  assign stOp_lane[1].scntl__dma__type0                     = scntl__sdp__lane1_type0                        ;
  assign stOp_lane[1].scntl__dma__num_of_types0             = scntl__sdp__lane1_num_of_types0                ;
  assign stOp_lane[2].scntl__dma__strm0_read_enable         = scntl__sdp__lane2_strm0_read_enable            ;
  assign stOp_lane[2].scntl__dma__strm0_write_enable        = scntl__sdp__lane2_strm0_write_enable           ;
  assign sdp__scntl__lane2_strm0_read_ready                 = stOp_lane[2].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane2_strm0_write_ready                = stOp_lane[2].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane2_strm0_read_complete              = stOp_lane[2].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane2_strm0_write_complete             = stOp_lane[2].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[2].scntl__dma__strm0_read_start_address  = scntl__sdp__lane2_strm0_read_start_address     ;
  assign stOp_lane[2].scntl__dma__strm0_write_start_address = scntl__sdp__lane2_strm0_write_start_address    ;
  assign stOp_lane[2].scntl__dma__type0                     = scntl__sdp__lane2_type0                        ;
  assign stOp_lane[2].scntl__dma__num_of_types0             = scntl__sdp__lane2_num_of_types0                ;
  assign stOp_lane[3].scntl__dma__strm0_read_enable         = scntl__sdp__lane3_strm0_read_enable            ;
  assign stOp_lane[3].scntl__dma__strm0_write_enable        = scntl__sdp__lane3_strm0_write_enable           ;
  assign sdp__scntl__lane3_strm0_read_ready                 = stOp_lane[3].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane3_strm0_write_ready                = stOp_lane[3].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane3_strm0_read_complete              = stOp_lane[3].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane3_strm0_write_complete             = stOp_lane[3].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[3].scntl__dma__strm0_read_start_address  = scntl__sdp__lane3_strm0_read_start_address     ;
  assign stOp_lane[3].scntl__dma__strm0_write_start_address = scntl__sdp__lane3_strm0_write_start_address    ;
  assign stOp_lane[3].scntl__dma__type0                     = scntl__sdp__lane3_type0                        ;
  assign stOp_lane[3].scntl__dma__num_of_types0             = scntl__sdp__lane3_num_of_types0                ;
  assign stOp_lane[4].scntl__dma__strm0_read_enable         = scntl__sdp__lane4_strm0_read_enable            ;
  assign stOp_lane[4].scntl__dma__strm0_write_enable        = scntl__sdp__lane4_strm0_write_enable           ;
  assign sdp__scntl__lane4_strm0_read_ready                 = stOp_lane[4].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane4_strm0_write_ready                = stOp_lane[4].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane4_strm0_read_complete              = stOp_lane[4].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane4_strm0_write_complete             = stOp_lane[4].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[4].scntl__dma__strm0_read_start_address  = scntl__sdp__lane4_strm0_read_start_address     ;
  assign stOp_lane[4].scntl__dma__strm0_write_start_address = scntl__sdp__lane4_strm0_write_start_address    ;
  assign stOp_lane[4].scntl__dma__type0                     = scntl__sdp__lane4_type0                        ;
  assign stOp_lane[4].scntl__dma__num_of_types0             = scntl__sdp__lane4_num_of_types0                ;
  assign stOp_lane[5].scntl__dma__strm0_read_enable         = scntl__sdp__lane5_strm0_read_enable            ;
  assign stOp_lane[5].scntl__dma__strm0_write_enable        = scntl__sdp__lane5_strm0_write_enable           ;
  assign sdp__scntl__lane5_strm0_read_ready                 = stOp_lane[5].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane5_strm0_write_ready                = stOp_lane[5].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane5_strm0_read_complete              = stOp_lane[5].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane5_strm0_write_complete             = stOp_lane[5].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[5].scntl__dma__strm0_read_start_address  = scntl__sdp__lane5_strm0_read_start_address     ;
  assign stOp_lane[5].scntl__dma__strm0_write_start_address = scntl__sdp__lane5_strm0_write_start_address    ;
  assign stOp_lane[5].scntl__dma__type0                     = scntl__sdp__lane5_type0                        ;
  assign stOp_lane[5].scntl__dma__num_of_types0             = scntl__sdp__lane5_num_of_types0                ;
  assign stOp_lane[6].scntl__dma__strm0_read_enable         = scntl__sdp__lane6_strm0_read_enable            ;
  assign stOp_lane[6].scntl__dma__strm0_write_enable        = scntl__sdp__lane6_strm0_write_enable           ;
  assign sdp__scntl__lane6_strm0_read_ready                 = stOp_lane[6].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane6_strm0_write_ready                = stOp_lane[6].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane6_strm0_read_complete              = stOp_lane[6].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane6_strm0_write_complete             = stOp_lane[6].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[6].scntl__dma__strm0_read_start_address  = scntl__sdp__lane6_strm0_read_start_address     ;
  assign stOp_lane[6].scntl__dma__strm0_write_start_address = scntl__sdp__lane6_strm0_write_start_address    ;
  assign stOp_lane[6].scntl__dma__type0                     = scntl__sdp__lane6_type0                        ;
  assign stOp_lane[6].scntl__dma__num_of_types0             = scntl__sdp__lane6_num_of_types0                ;
  assign stOp_lane[7].scntl__dma__strm0_read_enable         = scntl__sdp__lane7_strm0_read_enable            ;
  assign stOp_lane[7].scntl__dma__strm0_write_enable        = scntl__sdp__lane7_strm0_write_enable           ;
  assign sdp__scntl__lane7_strm0_read_ready                 = stOp_lane[7].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane7_strm0_write_ready                = stOp_lane[7].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane7_strm0_read_complete              = stOp_lane[7].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane7_strm0_write_complete             = stOp_lane[7].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[7].scntl__dma__strm0_read_start_address  = scntl__sdp__lane7_strm0_read_start_address     ;
  assign stOp_lane[7].scntl__dma__strm0_write_start_address = scntl__sdp__lane7_strm0_write_start_address    ;
  assign stOp_lane[7].scntl__dma__type0                     = scntl__sdp__lane7_type0                        ;
  assign stOp_lane[7].scntl__dma__num_of_types0             = scntl__sdp__lane7_num_of_types0                ;
  assign stOp_lane[8].scntl__dma__strm0_read_enable         = scntl__sdp__lane8_strm0_read_enable            ;
  assign stOp_lane[8].scntl__dma__strm0_write_enable        = scntl__sdp__lane8_strm0_write_enable           ;
  assign sdp__scntl__lane8_strm0_read_ready                 = stOp_lane[8].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane8_strm0_write_ready                = stOp_lane[8].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane8_strm0_read_complete              = stOp_lane[8].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane8_strm0_write_complete             = stOp_lane[8].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[8].scntl__dma__strm0_read_start_address  = scntl__sdp__lane8_strm0_read_start_address     ;
  assign stOp_lane[8].scntl__dma__strm0_write_start_address = scntl__sdp__lane8_strm0_write_start_address    ;
  assign stOp_lane[8].scntl__dma__type0                     = scntl__sdp__lane8_type0                        ;
  assign stOp_lane[8].scntl__dma__num_of_types0             = scntl__sdp__lane8_num_of_types0                ;
  assign stOp_lane[9].scntl__dma__strm0_read_enable         = scntl__sdp__lane9_strm0_read_enable            ;
  assign stOp_lane[9].scntl__dma__strm0_write_enable        = scntl__sdp__lane9_strm0_write_enable           ;
  assign sdp__scntl__lane9_strm0_read_ready                 = stOp_lane[9].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane9_strm0_write_ready                = stOp_lane[9].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane9_strm0_read_complete              = stOp_lane[9].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane9_strm0_write_complete             = stOp_lane[9].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[9].scntl__dma__strm0_read_start_address  = scntl__sdp__lane9_strm0_read_start_address     ;
  assign stOp_lane[9].scntl__dma__strm0_write_start_address = scntl__sdp__lane9_strm0_write_start_address    ;
  assign stOp_lane[9].scntl__dma__type0                     = scntl__sdp__lane9_type0                        ;
  assign stOp_lane[9].scntl__dma__num_of_types0             = scntl__sdp__lane9_num_of_types0                ;
  assign stOp_lane[10].scntl__dma__strm0_read_enable         = scntl__sdp__lane10_strm0_read_enable            ;
  assign stOp_lane[10].scntl__dma__strm0_write_enable        = scntl__sdp__lane10_strm0_write_enable           ;
  assign sdp__scntl__lane10_strm0_read_ready                 = stOp_lane[10].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane10_strm0_write_ready                = stOp_lane[10].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane10_strm0_read_complete              = stOp_lane[10].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane10_strm0_write_complete             = stOp_lane[10].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[10].scntl__dma__strm0_read_start_address  = scntl__sdp__lane10_strm0_read_start_address     ;
  assign stOp_lane[10].scntl__dma__strm0_write_start_address = scntl__sdp__lane10_strm0_write_start_address    ;
  assign stOp_lane[10].scntl__dma__type0                     = scntl__sdp__lane10_type0                        ;
  assign stOp_lane[10].scntl__dma__num_of_types0             = scntl__sdp__lane10_num_of_types0                ;
  assign stOp_lane[11].scntl__dma__strm0_read_enable         = scntl__sdp__lane11_strm0_read_enable            ;
  assign stOp_lane[11].scntl__dma__strm0_write_enable        = scntl__sdp__lane11_strm0_write_enable           ;
  assign sdp__scntl__lane11_strm0_read_ready                 = stOp_lane[11].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane11_strm0_write_ready                = stOp_lane[11].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane11_strm0_read_complete              = stOp_lane[11].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane11_strm0_write_complete             = stOp_lane[11].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[11].scntl__dma__strm0_read_start_address  = scntl__sdp__lane11_strm0_read_start_address     ;
  assign stOp_lane[11].scntl__dma__strm0_write_start_address = scntl__sdp__lane11_strm0_write_start_address    ;
  assign stOp_lane[11].scntl__dma__type0                     = scntl__sdp__lane11_type0                        ;
  assign stOp_lane[11].scntl__dma__num_of_types0             = scntl__sdp__lane11_num_of_types0                ;
  assign stOp_lane[12].scntl__dma__strm0_read_enable         = scntl__sdp__lane12_strm0_read_enable            ;
  assign stOp_lane[12].scntl__dma__strm0_write_enable        = scntl__sdp__lane12_strm0_write_enable           ;
  assign sdp__scntl__lane12_strm0_read_ready                 = stOp_lane[12].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane12_strm0_write_ready                = stOp_lane[12].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane12_strm0_read_complete              = stOp_lane[12].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane12_strm0_write_complete             = stOp_lane[12].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[12].scntl__dma__strm0_read_start_address  = scntl__sdp__lane12_strm0_read_start_address     ;
  assign stOp_lane[12].scntl__dma__strm0_write_start_address = scntl__sdp__lane12_strm0_write_start_address    ;
  assign stOp_lane[12].scntl__dma__type0                     = scntl__sdp__lane12_type0                        ;
  assign stOp_lane[12].scntl__dma__num_of_types0             = scntl__sdp__lane12_num_of_types0                ;
  assign stOp_lane[13].scntl__dma__strm0_read_enable         = scntl__sdp__lane13_strm0_read_enable            ;
  assign stOp_lane[13].scntl__dma__strm0_write_enable        = scntl__sdp__lane13_strm0_write_enable           ;
  assign sdp__scntl__lane13_strm0_read_ready                 = stOp_lane[13].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane13_strm0_write_ready                = stOp_lane[13].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane13_strm0_read_complete              = stOp_lane[13].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane13_strm0_write_complete             = stOp_lane[13].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[13].scntl__dma__strm0_read_start_address  = scntl__sdp__lane13_strm0_read_start_address     ;
  assign stOp_lane[13].scntl__dma__strm0_write_start_address = scntl__sdp__lane13_strm0_write_start_address    ;
  assign stOp_lane[13].scntl__dma__type0                     = scntl__sdp__lane13_type0                        ;
  assign stOp_lane[13].scntl__dma__num_of_types0             = scntl__sdp__lane13_num_of_types0                ;
  assign stOp_lane[14].scntl__dma__strm0_read_enable         = scntl__sdp__lane14_strm0_read_enable            ;
  assign stOp_lane[14].scntl__dma__strm0_write_enable        = scntl__sdp__lane14_strm0_write_enable           ;
  assign sdp__scntl__lane14_strm0_read_ready                 = stOp_lane[14].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane14_strm0_write_ready                = stOp_lane[14].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane14_strm0_read_complete              = stOp_lane[14].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane14_strm0_write_complete             = stOp_lane[14].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[14].scntl__dma__strm0_read_start_address  = scntl__sdp__lane14_strm0_read_start_address     ;
  assign stOp_lane[14].scntl__dma__strm0_write_start_address = scntl__sdp__lane14_strm0_write_start_address    ;
  assign stOp_lane[14].scntl__dma__type0                     = scntl__sdp__lane14_type0                        ;
  assign stOp_lane[14].scntl__dma__num_of_types0             = scntl__sdp__lane14_num_of_types0                ;
  assign stOp_lane[15].scntl__dma__strm0_read_enable         = scntl__sdp__lane15_strm0_read_enable            ;
  assign stOp_lane[15].scntl__dma__strm0_write_enable        = scntl__sdp__lane15_strm0_write_enable           ;
  assign sdp__scntl__lane15_strm0_read_ready                 = stOp_lane[15].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane15_strm0_write_ready                = stOp_lane[15].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane15_strm0_read_complete              = stOp_lane[15].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane15_strm0_write_complete             = stOp_lane[15].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[15].scntl__dma__strm0_read_start_address  = scntl__sdp__lane15_strm0_read_start_address     ;
  assign stOp_lane[15].scntl__dma__strm0_write_start_address = scntl__sdp__lane15_strm0_write_start_address    ;
  assign stOp_lane[15].scntl__dma__type0                     = scntl__sdp__lane15_type0                        ;
  assign stOp_lane[15].scntl__dma__num_of_types0             = scntl__sdp__lane15_num_of_types0                ;
  assign stOp_lane[16].scntl__dma__strm0_read_enable         = scntl__sdp__lane16_strm0_read_enable            ;
  assign stOp_lane[16].scntl__dma__strm0_write_enable        = scntl__sdp__lane16_strm0_write_enable           ;
  assign sdp__scntl__lane16_strm0_read_ready                 = stOp_lane[16].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane16_strm0_write_ready                = stOp_lane[16].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane16_strm0_read_complete              = stOp_lane[16].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane16_strm0_write_complete             = stOp_lane[16].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[16].scntl__dma__strm0_read_start_address  = scntl__sdp__lane16_strm0_read_start_address     ;
  assign stOp_lane[16].scntl__dma__strm0_write_start_address = scntl__sdp__lane16_strm0_write_start_address    ;
  assign stOp_lane[16].scntl__dma__type0                     = scntl__sdp__lane16_type0                        ;
  assign stOp_lane[16].scntl__dma__num_of_types0             = scntl__sdp__lane16_num_of_types0                ;
  assign stOp_lane[17].scntl__dma__strm0_read_enable         = scntl__sdp__lane17_strm0_read_enable            ;
  assign stOp_lane[17].scntl__dma__strm0_write_enable        = scntl__sdp__lane17_strm0_write_enable           ;
  assign sdp__scntl__lane17_strm0_read_ready                 = stOp_lane[17].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane17_strm0_write_ready                = stOp_lane[17].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane17_strm0_read_complete              = stOp_lane[17].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane17_strm0_write_complete             = stOp_lane[17].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[17].scntl__dma__strm0_read_start_address  = scntl__sdp__lane17_strm0_read_start_address     ;
  assign stOp_lane[17].scntl__dma__strm0_write_start_address = scntl__sdp__lane17_strm0_write_start_address    ;
  assign stOp_lane[17].scntl__dma__type0                     = scntl__sdp__lane17_type0                        ;
  assign stOp_lane[17].scntl__dma__num_of_types0             = scntl__sdp__lane17_num_of_types0                ;
  assign stOp_lane[18].scntl__dma__strm0_read_enable         = scntl__sdp__lane18_strm0_read_enable            ;
  assign stOp_lane[18].scntl__dma__strm0_write_enable        = scntl__sdp__lane18_strm0_write_enable           ;
  assign sdp__scntl__lane18_strm0_read_ready                 = stOp_lane[18].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane18_strm0_write_ready                = stOp_lane[18].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane18_strm0_read_complete              = stOp_lane[18].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane18_strm0_write_complete             = stOp_lane[18].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[18].scntl__dma__strm0_read_start_address  = scntl__sdp__lane18_strm0_read_start_address     ;
  assign stOp_lane[18].scntl__dma__strm0_write_start_address = scntl__sdp__lane18_strm0_write_start_address    ;
  assign stOp_lane[18].scntl__dma__type0                     = scntl__sdp__lane18_type0                        ;
  assign stOp_lane[18].scntl__dma__num_of_types0             = scntl__sdp__lane18_num_of_types0                ;
  assign stOp_lane[19].scntl__dma__strm0_read_enable         = scntl__sdp__lane19_strm0_read_enable            ;
  assign stOp_lane[19].scntl__dma__strm0_write_enable        = scntl__sdp__lane19_strm0_write_enable           ;
  assign sdp__scntl__lane19_strm0_read_ready                 = stOp_lane[19].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane19_strm0_write_ready                = stOp_lane[19].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane19_strm0_read_complete              = stOp_lane[19].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane19_strm0_write_complete             = stOp_lane[19].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[19].scntl__dma__strm0_read_start_address  = scntl__sdp__lane19_strm0_read_start_address     ;
  assign stOp_lane[19].scntl__dma__strm0_write_start_address = scntl__sdp__lane19_strm0_write_start_address    ;
  assign stOp_lane[19].scntl__dma__type0                     = scntl__sdp__lane19_type0                        ;
  assign stOp_lane[19].scntl__dma__num_of_types0             = scntl__sdp__lane19_num_of_types0                ;
  assign stOp_lane[20].scntl__dma__strm0_read_enable         = scntl__sdp__lane20_strm0_read_enable            ;
  assign stOp_lane[20].scntl__dma__strm0_write_enable        = scntl__sdp__lane20_strm0_write_enable           ;
  assign sdp__scntl__lane20_strm0_read_ready                 = stOp_lane[20].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane20_strm0_write_ready                = stOp_lane[20].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane20_strm0_read_complete              = stOp_lane[20].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane20_strm0_write_complete             = stOp_lane[20].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[20].scntl__dma__strm0_read_start_address  = scntl__sdp__lane20_strm0_read_start_address     ;
  assign stOp_lane[20].scntl__dma__strm0_write_start_address = scntl__sdp__lane20_strm0_write_start_address    ;
  assign stOp_lane[20].scntl__dma__type0                     = scntl__sdp__lane20_type0                        ;
  assign stOp_lane[20].scntl__dma__num_of_types0             = scntl__sdp__lane20_num_of_types0                ;
  assign stOp_lane[21].scntl__dma__strm0_read_enable         = scntl__sdp__lane21_strm0_read_enable            ;
  assign stOp_lane[21].scntl__dma__strm0_write_enable        = scntl__sdp__lane21_strm0_write_enable           ;
  assign sdp__scntl__lane21_strm0_read_ready                 = stOp_lane[21].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane21_strm0_write_ready                = stOp_lane[21].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane21_strm0_read_complete              = stOp_lane[21].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane21_strm0_write_complete             = stOp_lane[21].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[21].scntl__dma__strm0_read_start_address  = scntl__sdp__lane21_strm0_read_start_address     ;
  assign stOp_lane[21].scntl__dma__strm0_write_start_address = scntl__sdp__lane21_strm0_write_start_address    ;
  assign stOp_lane[21].scntl__dma__type0                     = scntl__sdp__lane21_type0                        ;
  assign stOp_lane[21].scntl__dma__num_of_types0             = scntl__sdp__lane21_num_of_types0                ;
  assign stOp_lane[22].scntl__dma__strm0_read_enable         = scntl__sdp__lane22_strm0_read_enable            ;
  assign stOp_lane[22].scntl__dma__strm0_write_enable        = scntl__sdp__lane22_strm0_write_enable           ;
  assign sdp__scntl__lane22_strm0_read_ready                 = stOp_lane[22].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane22_strm0_write_ready                = stOp_lane[22].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane22_strm0_read_complete              = stOp_lane[22].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane22_strm0_write_complete             = stOp_lane[22].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[22].scntl__dma__strm0_read_start_address  = scntl__sdp__lane22_strm0_read_start_address     ;
  assign stOp_lane[22].scntl__dma__strm0_write_start_address = scntl__sdp__lane22_strm0_write_start_address    ;
  assign stOp_lane[22].scntl__dma__type0                     = scntl__sdp__lane22_type0                        ;
  assign stOp_lane[22].scntl__dma__num_of_types0             = scntl__sdp__lane22_num_of_types0                ;
  assign stOp_lane[23].scntl__dma__strm0_read_enable         = scntl__sdp__lane23_strm0_read_enable            ;
  assign stOp_lane[23].scntl__dma__strm0_write_enable        = scntl__sdp__lane23_strm0_write_enable           ;
  assign sdp__scntl__lane23_strm0_read_ready                 = stOp_lane[23].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane23_strm0_write_ready                = stOp_lane[23].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane23_strm0_read_complete              = stOp_lane[23].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane23_strm0_write_complete             = stOp_lane[23].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[23].scntl__dma__strm0_read_start_address  = scntl__sdp__lane23_strm0_read_start_address     ;
  assign stOp_lane[23].scntl__dma__strm0_write_start_address = scntl__sdp__lane23_strm0_write_start_address    ;
  assign stOp_lane[23].scntl__dma__type0                     = scntl__sdp__lane23_type0                        ;
  assign stOp_lane[23].scntl__dma__num_of_types0             = scntl__sdp__lane23_num_of_types0                ;
  assign stOp_lane[24].scntl__dma__strm0_read_enable         = scntl__sdp__lane24_strm0_read_enable            ;
  assign stOp_lane[24].scntl__dma__strm0_write_enable        = scntl__sdp__lane24_strm0_write_enable           ;
  assign sdp__scntl__lane24_strm0_read_ready                 = stOp_lane[24].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane24_strm0_write_ready                = stOp_lane[24].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane24_strm0_read_complete              = stOp_lane[24].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane24_strm0_write_complete             = stOp_lane[24].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[24].scntl__dma__strm0_read_start_address  = scntl__sdp__lane24_strm0_read_start_address     ;
  assign stOp_lane[24].scntl__dma__strm0_write_start_address = scntl__sdp__lane24_strm0_write_start_address    ;
  assign stOp_lane[24].scntl__dma__type0                     = scntl__sdp__lane24_type0                        ;
  assign stOp_lane[24].scntl__dma__num_of_types0             = scntl__sdp__lane24_num_of_types0                ;
  assign stOp_lane[25].scntl__dma__strm0_read_enable         = scntl__sdp__lane25_strm0_read_enable            ;
  assign stOp_lane[25].scntl__dma__strm0_write_enable        = scntl__sdp__lane25_strm0_write_enable           ;
  assign sdp__scntl__lane25_strm0_read_ready                 = stOp_lane[25].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane25_strm0_write_ready                = stOp_lane[25].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane25_strm0_read_complete              = stOp_lane[25].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane25_strm0_write_complete             = stOp_lane[25].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[25].scntl__dma__strm0_read_start_address  = scntl__sdp__lane25_strm0_read_start_address     ;
  assign stOp_lane[25].scntl__dma__strm0_write_start_address = scntl__sdp__lane25_strm0_write_start_address    ;
  assign stOp_lane[25].scntl__dma__type0                     = scntl__sdp__lane25_type0                        ;
  assign stOp_lane[25].scntl__dma__num_of_types0             = scntl__sdp__lane25_num_of_types0                ;
  assign stOp_lane[26].scntl__dma__strm0_read_enable         = scntl__sdp__lane26_strm0_read_enable            ;
  assign stOp_lane[26].scntl__dma__strm0_write_enable        = scntl__sdp__lane26_strm0_write_enable           ;
  assign sdp__scntl__lane26_strm0_read_ready                 = stOp_lane[26].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane26_strm0_write_ready                = stOp_lane[26].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane26_strm0_read_complete              = stOp_lane[26].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane26_strm0_write_complete             = stOp_lane[26].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[26].scntl__dma__strm0_read_start_address  = scntl__sdp__lane26_strm0_read_start_address     ;
  assign stOp_lane[26].scntl__dma__strm0_write_start_address = scntl__sdp__lane26_strm0_write_start_address    ;
  assign stOp_lane[26].scntl__dma__type0                     = scntl__sdp__lane26_type0                        ;
  assign stOp_lane[26].scntl__dma__num_of_types0             = scntl__sdp__lane26_num_of_types0                ;
  assign stOp_lane[27].scntl__dma__strm0_read_enable         = scntl__sdp__lane27_strm0_read_enable            ;
  assign stOp_lane[27].scntl__dma__strm0_write_enable        = scntl__sdp__lane27_strm0_write_enable           ;
  assign sdp__scntl__lane27_strm0_read_ready                 = stOp_lane[27].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane27_strm0_write_ready                = stOp_lane[27].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane27_strm0_read_complete              = stOp_lane[27].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane27_strm0_write_complete             = stOp_lane[27].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[27].scntl__dma__strm0_read_start_address  = scntl__sdp__lane27_strm0_read_start_address     ;
  assign stOp_lane[27].scntl__dma__strm0_write_start_address = scntl__sdp__lane27_strm0_write_start_address    ;
  assign stOp_lane[27].scntl__dma__type0                     = scntl__sdp__lane27_type0                        ;
  assign stOp_lane[27].scntl__dma__num_of_types0             = scntl__sdp__lane27_num_of_types0                ;
  assign stOp_lane[28].scntl__dma__strm0_read_enable         = scntl__sdp__lane28_strm0_read_enable            ;
  assign stOp_lane[28].scntl__dma__strm0_write_enable        = scntl__sdp__lane28_strm0_write_enable           ;
  assign sdp__scntl__lane28_strm0_read_ready                 = stOp_lane[28].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane28_strm0_write_ready                = stOp_lane[28].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane28_strm0_read_complete              = stOp_lane[28].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane28_strm0_write_complete             = stOp_lane[28].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[28].scntl__dma__strm0_read_start_address  = scntl__sdp__lane28_strm0_read_start_address     ;
  assign stOp_lane[28].scntl__dma__strm0_write_start_address = scntl__sdp__lane28_strm0_write_start_address    ;
  assign stOp_lane[28].scntl__dma__type0                     = scntl__sdp__lane28_type0                        ;
  assign stOp_lane[28].scntl__dma__num_of_types0             = scntl__sdp__lane28_num_of_types0                ;
  assign stOp_lane[29].scntl__dma__strm0_read_enable         = scntl__sdp__lane29_strm0_read_enable            ;
  assign stOp_lane[29].scntl__dma__strm0_write_enable        = scntl__sdp__lane29_strm0_write_enable           ;
  assign sdp__scntl__lane29_strm0_read_ready                 = stOp_lane[29].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane29_strm0_write_ready                = stOp_lane[29].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane29_strm0_read_complete              = stOp_lane[29].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane29_strm0_write_complete             = stOp_lane[29].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[29].scntl__dma__strm0_read_start_address  = scntl__sdp__lane29_strm0_read_start_address     ;
  assign stOp_lane[29].scntl__dma__strm0_write_start_address = scntl__sdp__lane29_strm0_write_start_address    ;
  assign stOp_lane[29].scntl__dma__type0                     = scntl__sdp__lane29_type0                        ;
  assign stOp_lane[29].scntl__dma__num_of_types0             = scntl__sdp__lane29_num_of_types0                ;
  assign stOp_lane[30].scntl__dma__strm0_read_enable         = scntl__sdp__lane30_strm0_read_enable            ;
  assign stOp_lane[30].scntl__dma__strm0_write_enable        = scntl__sdp__lane30_strm0_write_enable           ;
  assign sdp__scntl__lane30_strm0_read_ready                 = stOp_lane[30].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane30_strm0_write_ready                = stOp_lane[30].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane30_strm0_read_complete              = stOp_lane[30].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane30_strm0_write_complete             = stOp_lane[30].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[30].scntl__dma__strm0_read_start_address  = scntl__sdp__lane30_strm0_read_start_address     ;
  assign stOp_lane[30].scntl__dma__strm0_write_start_address = scntl__sdp__lane30_strm0_write_start_address    ;
  assign stOp_lane[30].scntl__dma__type0                     = scntl__sdp__lane30_type0                        ;
  assign stOp_lane[30].scntl__dma__num_of_types0             = scntl__sdp__lane30_num_of_types0                ;
  assign stOp_lane[31].scntl__dma__strm0_read_enable         = scntl__sdp__lane31_strm0_read_enable            ;
  assign stOp_lane[31].scntl__dma__strm0_write_enable        = scntl__sdp__lane31_strm0_write_enable           ;
  assign sdp__scntl__lane31_strm0_read_ready                 = stOp_lane[31].dma__scntl__strm0_read_ready      ;
  assign sdp__scntl__lane31_strm0_write_ready                = stOp_lane[31].dma__scntl__strm0_write_ready     ;
  assign sdp__scntl__lane31_strm0_read_complete              = stOp_lane[31].dma__scntl__strm0_read_complete   ;
  assign sdp__scntl__lane31_strm0_write_complete             = stOp_lane[31].dma__scntl__strm0_write_complete  ;
  assign stOp_lane[31].scntl__dma__strm0_read_start_address  = scntl__sdp__lane31_strm0_read_start_address     ;
  assign stOp_lane[31].scntl__dma__strm0_write_start_address = scntl__sdp__lane31_strm0_write_start_address    ;
  assign stOp_lane[31].scntl__dma__type0                     = scntl__sdp__lane31_type0                        ;
  assign stOp_lane[31].scntl__dma__num_of_types0             = scntl__sdp__lane31_num_of_types0                ;
