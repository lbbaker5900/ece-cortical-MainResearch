
  assign  mgr0__std__oob_cntl                       =  mgr_inst[0].mgr__std__oob_cntl       ;
  assign  mgr0__std__oob_valid                      =  mgr_inst[0].mgr__std__oob_valid      ;
  assign  mgr_inst[0].std__mgr__oob_ready           =  std__mgr0__oob_ready                 ;
  assign  mgr0__std__oob_type                       =  mgr_inst[0].mgr__std__oob_type       ;
  assign  mgr0__std__oob_data                       =  mgr_inst[0].mgr__std__oob_data       ;

  assign  mgr1__std__oob_cntl                       =  mgr_inst[1].mgr__std__oob_cntl       ;
  assign  mgr1__std__oob_valid                      =  mgr_inst[1].mgr__std__oob_valid      ;
  assign  mgr_inst[1].std__mgr__oob_ready           =  std__mgr1__oob_ready                 ;
  assign  mgr1__std__oob_type                       =  mgr_inst[1].mgr__std__oob_type       ;
  assign  mgr1__std__oob_data                       =  mgr_inst[1].mgr__std__oob_data       ;

  assign  mgr2__std__oob_cntl                       =  mgr_inst[2].mgr__std__oob_cntl       ;
  assign  mgr2__std__oob_valid                      =  mgr_inst[2].mgr__std__oob_valid      ;
  assign  mgr_inst[2].std__mgr__oob_ready           =  std__mgr2__oob_ready                 ;
  assign  mgr2__std__oob_type                       =  mgr_inst[2].mgr__std__oob_type       ;
  assign  mgr2__std__oob_data                       =  mgr_inst[2].mgr__std__oob_data       ;

  assign  mgr3__std__oob_cntl                       =  mgr_inst[3].mgr__std__oob_cntl       ;
  assign  mgr3__std__oob_valid                      =  mgr_inst[3].mgr__std__oob_valid      ;
  assign  mgr_inst[3].std__mgr__oob_ready           =  std__mgr3__oob_ready                 ;
  assign  mgr3__std__oob_type                       =  mgr_inst[3].mgr__std__oob_type       ;
  assign  mgr3__std__oob_data                       =  mgr_inst[3].mgr__std__oob_data       ;

