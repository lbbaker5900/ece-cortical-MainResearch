
    .reg__scntl__ready [0]   ( reg__scntl__lane0_ready  ) ,
    .scntl__reg__valid [0]   ( scntl__reg__lane0_valid  ) ,
    .scntl__reg__data  [0]   ( scntl__reg__lane0_data   ) ,

    .reg__scntl__ready [1]   ( reg__scntl__lane1_ready  ) ,
    .scntl__reg__valid [1]   ( scntl__reg__lane1_valid  ) ,
    .scntl__reg__data  [1]   ( scntl__reg__lane1_data   ) ,

    .reg__scntl__ready [2]   ( reg__scntl__lane2_ready  ) ,
    .scntl__reg__valid [2]   ( scntl__reg__lane2_valid  ) ,
    .scntl__reg__data  [2]   ( scntl__reg__lane2_data   ) ,

    .reg__scntl__ready [3]   ( reg__scntl__lane3_ready  ) ,
    .scntl__reg__valid [3]   ( scntl__reg__lane3_valid  ) ,
    .scntl__reg__data  [3]   ( scntl__reg__lane3_data   ) ,

    .reg__scntl__ready [4]   ( reg__scntl__lane4_ready  ) ,
    .scntl__reg__valid [4]   ( scntl__reg__lane4_valid  ) ,
    .scntl__reg__data  [4]   ( scntl__reg__lane4_data   ) ,

    .reg__scntl__ready [5]   ( reg__scntl__lane5_ready  ) ,
    .scntl__reg__valid [5]   ( scntl__reg__lane5_valid  ) ,
    .scntl__reg__data  [5]   ( scntl__reg__lane5_data   ) ,

    .reg__scntl__ready [6]   ( reg__scntl__lane6_ready  ) ,
    .scntl__reg__valid [6]   ( scntl__reg__lane6_valid  ) ,
    .scntl__reg__data  [6]   ( scntl__reg__lane6_data   ) ,

    .reg__scntl__ready [7]   ( reg__scntl__lane7_ready  ) ,
    .scntl__reg__valid [7]   ( scntl__reg__lane7_valid  ) ,
    .scntl__reg__data  [7]   ( scntl__reg__lane7_data   ) ,

    .reg__scntl__ready [8]   ( reg__scntl__lane8_ready  ) ,
    .scntl__reg__valid [8]   ( scntl__reg__lane8_valid  ) ,
    .scntl__reg__data  [8]   ( scntl__reg__lane8_data   ) ,

    .reg__scntl__ready [9]   ( reg__scntl__lane9_ready  ) ,
    .scntl__reg__valid [9]   ( scntl__reg__lane9_valid  ) ,
    .scntl__reg__data  [9]   ( scntl__reg__lane9_data   ) ,

    .reg__scntl__ready [10]   ( reg__scntl__lane10_ready  ) ,
    .scntl__reg__valid [10]   ( scntl__reg__lane10_valid  ) ,
    .scntl__reg__data  [10]   ( scntl__reg__lane10_data   ) ,

    .reg__scntl__ready [11]   ( reg__scntl__lane11_ready  ) ,
    .scntl__reg__valid [11]   ( scntl__reg__lane11_valid  ) ,
    .scntl__reg__data  [11]   ( scntl__reg__lane11_data   ) ,

    .reg__scntl__ready [12]   ( reg__scntl__lane12_ready  ) ,
    .scntl__reg__valid [12]   ( scntl__reg__lane12_valid  ) ,
    .scntl__reg__data  [12]   ( scntl__reg__lane12_data   ) ,

    .reg__scntl__ready [13]   ( reg__scntl__lane13_ready  ) ,
    .scntl__reg__valid [13]   ( scntl__reg__lane13_valid  ) ,
    .scntl__reg__data  [13]   ( scntl__reg__lane13_data   ) ,

    .reg__scntl__ready [14]   ( reg__scntl__lane14_ready  ) ,
    .scntl__reg__valid [14]   ( scntl__reg__lane14_valid  ) ,
    .scntl__reg__data  [14]   ( scntl__reg__lane14_data   ) ,

    .reg__scntl__ready [15]   ( reg__scntl__lane15_ready  ) ,
    .scntl__reg__valid [15]   ( scntl__reg__lane15_valid  ) ,
    .scntl__reg__data  [15]   ( scntl__reg__lane15_data   ) ,

    .reg__scntl__ready [16]   ( reg__scntl__lane16_ready  ) ,
    .scntl__reg__valid [16]   ( scntl__reg__lane16_valid  ) ,
    .scntl__reg__data  [16]   ( scntl__reg__lane16_data   ) ,

    .reg__scntl__ready [17]   ( reg__scntl__lane17_ready  ) ,
    .scntl__reg__valid [17]   ( scntl__reg__lane17_valid  ) ,
    .scntl__reg__data  [17]   ( scntl__reg__lane17_data   ) ,

    .reg__scntl__ready [18]   ( reg__scntl__lane18_ready  ) ,
    .scntl__reg__valid [18]   ( scntl__reg__lane18_valid  ) ,
    .scntl__reg__data  [18]   ( scntl__reg__lane18_data   ) ,

    .reg__scntl__ready [19]   ( reg__scntl__lane19_ready  ) ,
    .scntl__reg__valid [19]   ( scntl__reg__lane19_valid  ) ,
    .scntl__reg__data  [19]   ( scntl__reg__lane19_data   ) ,

    .reg__scntl__ready [20]   ( reg__scntl__lane20_ready  ) ,
    .scntl__reg__valid [20]   ( scntl__reg__lane20_valid  ) ,
    .scntl__reg__data  [20]   ( scntl__reg__lane20_data   ) ,

    .reg__scntl__ready [21]   ( reg__scntl__lane21_ready  ) ,
    .scntl__reg__valid [21]   ( scntl__reg__lane21_valid  ) ,
    .scntl__reg__data  [21]   ( scntl__reg__lane21_data   ) ,

    .reg__scntl__ready [22]   ( reg__scntl__lane22_ready  ) ,
    .scntl__reg__valid [22]   ( scntl__reg__lane22_valid  ) ,
    .scntl__reg__data  [22]   ( scntl__reg__lane22_data   ) ,

    .reg__scntl__ready [23]   ( reg__scntl__lane23_ready  ) ,
    .scntl__reg__valid [23]   ( scntl__reg__lane23_valid  ) ,
    .scntl__reg__data  [23]   ( scntl__reg__lane23_data   ) ,

    .reg__scntl__ready [24]   ( reg__scntl__lane24_ready  ) ,
    .scntl__reg__valid [24]   ( scntl__reg__lane24_valid  ) ,
    .scntl__reg__data  [24]   ( scntl__reg__lane24_data   ) ,

    .reg__scntl__ready [25]   ( reg__scntl__lane25_ready  ) ,
    .scntl__reg__valid [25]   ( scntl__reg__lane25_valid  ) ,
    .scntl__reg__data  [25]   ( scntl__reg__lane25_data   ) ,

    .reg__scntl__ready [26]   ( reg__scntl__lane26_ready  ) ,
    .scntl__reg__valid [26]   ( scntl__reg__lane26_valid  ) ,
    .scntl__reg__data  [26]   ( scntl__reg__lane26_data   ) ,

    .reg__scntl__ready [27]   ( reg__scntl__lane27_ready  ) ,
    .scntl__reg__valid [27]   ( scntl__reg__lane27_valid  ) ,
    .scntl__reg__data  [27]   ( scntl__reg__lane27_data   ) ,

    .reg__scntl__ready [28]   ( reg__scntl__lane28_ready  ) ,
    .scntl__reg__valid [28]   ( scntl__reg__lane28_valid  ) ,
    .scntl__reg__data  [28]   ( scntl__reg__lane28_data   ) ,

    .reg__scntl__ready [29]   ( reg__scntl__lane29_ready  ) ,
    .scntl__reg__valid [29]   ( scntl__reg__lane29_valid  ) ,
    .scntl__reg__data  [29]   ( scntl__reg__lane29_data   ) ,

    .reg__scntl__ready [30]   ( reg__scntl__lane30_ready  ) ,
    .scntl__reg__valid [30]   ( scntl__reg__lane30_valid  ) ,
    .scntl__reg__data  [30]   ( scntl__reg__lane30_data   ) ,

    .reg__scntl__ready [31]   ( reg__scntl__lane31_ready  ) ,
    .scntl__reg__valid [31]   ( scntl__reg__lane31_valid  ) ,
    .scntl__reg__data  [31]   ( scntl__reg__lane31_data   ) ,

