
  // General control and status                                                 
  wire                                        mgr0__sys__allSynchronized     ;
  wire                                        sys__mgr0__thisSynchronized    ;
  wire                                        sys__mgr0__ready               ;
  wire                                        sys__mgr0__complete            ;

  // General control and status                                                 
  wire                                        mgr1__sys__allSynchronized     ;
  wire                                        sys__mgr1__thisSynchronized    ;
  wire                                        sys__mgr1__ready               ;
  wire                                        sys__mgr1__complete            ;

  // General control and status                                                 
  wire                                        mgr2__sys__allSynchronized     ;
  wire                                        sys__mgr2__thisSynchronized    ;
  wire                                        sys__mgr2__ready               ;
  wire                                        sys__mgr2__complete            ;

  // General control and status                                                 
  wire                                        mgr3__sys__allSynchronized     ;
  wire                                        sys__mgr3__thisSynchronized    ;
  wire                                        sys__mgr3__ready               ;
  wire                                        sys__mgr3__complete            ;
