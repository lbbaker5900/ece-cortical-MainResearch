
  output                                   reg__sdp__lane0_ready    ;
  input                                    sdp__reg__lane0_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane0_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane0_data     ;

  output                                   reg__sdp__lane1_ready    ;
  input                                    sdp__reg__lane1_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane1_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane1_data     ;

  output                                   reg__sdp__lane2_ready    ;
  input                                    sdp__reg__lane2_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane2_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane2_data     ;

  output                                   reg__sdp__lane3_ready    ;
  input                                    sdp__reg__lane3_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane3_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane3_data     ;

  output                                   reg__sdp__lane4_ready    ;
  input                                    sdp__reg__lane4_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane4_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane4_data     ;

  output                                   reg__sdp__lane5_ready    ;
  input                                    sdp__reg__lane5_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane5_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane5_data     ;

  output                                   reg__sdp__lane6_ready    ;
  input                                    sdp__reg__lane6_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane6_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane6_data     ;

  output                                   reg__sdp__lane7_ready    ;
  input                                    sdp__reg__lane7_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane7_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane7_data     ;

  output                                   reg__sdp__lane8_ready    ;
  input                                    sdp__reg__lane8_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane8_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane8_data     ;

  output                                   reg__sdp__lane9_ready    ;
  input                                    sdp__reg__lane9_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane9_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane9_data     ;

  output                                   reg__sdp__lane10_ready    ;
  input                                    sdp__reg__lane10_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane10_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane10_data     ;

  output                                   reg__sdp__lane11_ready    ;
  input                                    sdp__reg__lane11_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane11_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane11_data     ;

  output                                   reg__sdp__lane12_ready    ;
  input                                    sdp__reg__lane12_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane12_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane12_data     ;

  output                                   reg__sdp__lane13_ready    ;
  input                                    sdp__reg__lane13_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane13_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane13_data     ;

  output                                   reg__sdp__lane14_ready    ;
  input                                    sdp__reg__lane14_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane14_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane14_data     ;

  output                                   reg__sdp__lane15_ready    ;
  input                                    sdp__reg__lane15_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane15_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane15_data     ;

  output                                   reg__sdp__lane16_ready    ;
  input                                    sdp__reg__lane16_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane16_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane16_data     ;

  output                                   reg__sdp__lane17_ready    ;
  input                                    sdp__reg__lane17_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane17_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane17_data     ;

  output                                   reg__sdp__lane18_ready    ;
  input                                    sdp__reg__lane18_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane18_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane18_data     ;

  output                                   reg__sdp__lane19_ready    ;
  input                                    sdp__reg__lane19_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane19_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane19_data     ;

  output                                   reg__sdp__lane20_ready    ;
  input                                    sdp__reg__lane20_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane20_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane20_data     ;

  output                                   reg__sdp__lane21_ready    ;
  input                                    sdp__reg__lane21_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane21_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane21_data     ;

  output                                   reg__sdp__lane22_ready    ;
  input                                    sdp__reg__lane22_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane22_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane22_data     ;

  output                                   reg__sdp__lane23_ready    ;
  input                                    sdp__reg__lane23_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane23_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane23_data     ;

  output                                   reg__sdp__lane24_ready    ;
  input                                    sdp__reg__lane24_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane24_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane24_data     ;

  output                                   reg__sdp__lane25_ready    ;
  input                                    sdp__reg__lane25_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane25_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane25_data     ;

  output                                   reg__sdp__lane26_ready    ;
  input                                    sdp__reg__lane26_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane26_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane26_data     ;

  output                                   reg__sdp__lane27_ready    ;
  input                                    sdp__reg__lane27_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane27_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane27_data     ;

  output                                   reg__sdp__lane28_ready    ;
  input                                    sdp__reg__lane28_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane28_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane28_data     ;

  output                                   reg__sdp__lane29_ready    ;
  input                                    sdp__reg__lane29_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane29_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane29_data     ;

  output                                   reg__sdp__lane30_ready    ;
  input                                    sdp__reg__lane30_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane30_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane30_data     ;

  output                                   reg__sdp__lane31_ready    ;
  input                                    sdp__reg__lane31_valid    ;
  input   [`COMMON_STD_INTF_CNTL_RANGE  ]  sdp__reg__lane31_cntl     ;
  input   [`STREAMING_OP_RESULT_RANGE   ]  sdp__reg__lane31_data     ;

