`define MGR_NOC_CONT_MGR0_PORT0_DESTINATION_MGR_BITMASK  'b10_10
`define MGR_NOC_CONT_MGR0_PORT1_DESTINATION_MGR_BITMASK  'b01_00
`define MGR_NOC_CONT_MGR0_PORT2_DESTINATION_MGR_BITMASK  'd0
`define MGR_NOC_CONT_MGR0_PORT3_DESTINATION_MGR_BITMASK  'd0
`define MGR_NOC_CONT_MGR1_PORT0_DESTINATION_MGR_BITMASK  'b10_00
`define MGR_NOC_CONT_MGR1_PORT1_DESTINATION_MGR_BITMASK  'b01_01
`define MGR_NOC_CONT_MGR1_PORT2_DESTINATION_MGR_BITMASK  'd0
`define MGR_NOC_CONT_MGR1_PORT3_DESTINATION_MGR_BITMASK  'd0
`define MGR_NOC_CONT_MGR2_PORT0_DESTINATION_MGR_BITMASK  'b00_11
`define MGR_NOC_CONT_MGR2_PORT1_DESTINATION_MGR_BITMASK  'b10_00
`define MGR_NOC_CONT_MGR2_PORT2_DESTINATION_MGR_BITMASK  'd0
`define MGR_NOC_CONT_MGR2_PORT3_DESTINATION_MGR_BITMASK  'd0
`define MGR_NOC_CONT_MGR3_PORT0_DESTINATION_MGR_BITMASK  'b00_11
`define MGR_NOC_CONT_MGR3_PORT1_DESTINATION_MGR_BITMASK  'b01_00
`define MGR_NOC_CONT_MGR3_PORT2_DESTINATION_MGR_BITMASK  'd0
`define MGR_NOC_CONT_MGR3_PORT3_DESTINATION_MGR_BITMASK  'd0
