
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[0] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[0] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[0].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[0].Id[1]  =  0      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[0].put(sys_operation_lane[0])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[0].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[0];                                                                                                                
            join_none                                                                                                                             
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[1] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[1] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[1].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[1].Id[1]  =  1      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[1].put(sys_operation_lane[1])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[1].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[1];                                                                                                                
            join_none                                                                                                                             
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[2] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[2] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[2].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[2].Id[1]  =  2      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[2].put(sys_operation_lane[2])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[2].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[2];                                                                                                                
            join_none                                                                                                                             
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[3] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[3] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[3].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[3].Id[1]  =  3      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[3].put(sys_operation_lane[3])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[3].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[3];                                                                                                                
            join_none                                                                                                                             
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[4] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[4] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[4].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[4].Id[1]  =  4      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[4].put(sys_operation_lane[4])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[4].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[4];                                                                                                                
            join_none                                                                                                                             
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[5] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[5] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[5].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[5].Id[1]  =  5      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[5].put(sys_operation_lane[5])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[5].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[5];                                                                                                                
            join_none                                                                                                                             
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[6] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[6] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[6].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[6].Id[1]  =  6      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[6].put(sys_operation_lane[6])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[6].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[6];                                                                                                                
            join_none                                                                                                                             
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[7] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[7] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[7].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[7].Id[1]  =  7      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[7].put(sys_operation_lane[7])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[7].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[7];                                                                                                                
            join_none                                                                                                                             
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[8] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[8] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[8].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[8].Id[1]  =  8      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[8].put(sys_operation_lane[8])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[8].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[8];                                                                                                                
            join_none                                                                                                                             
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[9] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[9] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[9].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[9].Id[1]  =  9      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[9].put(sys_operation_lane[9])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[9].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[9];                                                                                                                
            join_none                                                                                                                             
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[10] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[10] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[10].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[10].Id[1]  =  10      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[10].put(sys_operation_lane[10])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[10].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[10];                                                                                                                
            join_none                                                                                                                             
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[11] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[11] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[11].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[11].Id[1]  =  11      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[11].put(sys_operation_lane[11])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[11].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[11];                                                                                                                
            join_none                                                                                                                             
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[12] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[12] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[12].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[12].Id[1]  =  12      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[12].put(sys_operation_lane[12])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[12].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[12];                                                                                                                
            join_none                                                                                                                             
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[13] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[13] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[13].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[13].Id[1]  =  13      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[13].put(sys_operation_lane[13])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[13].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[13];                                                                                                                
            join_none                                                                                                                             
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[14] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[14] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[14].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[14].Id[1]  =  14      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[14].put(sys_operation_lane[14])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[14].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[14];                                                                                                                
            join_none                                                                                                                             
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[15] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[15] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[15].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[15].Id[1]  =  15      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[15].put(sys_operation_lane[15])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[15].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[15];                                                                                                                
            join_none                                                                                                                             
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[16] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[16] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[16].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[16].Id[1]  =  16      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[16].put(sys_operation_lane[16])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[16].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[16];                                                                                                                
            join_none                                                                                                                             
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[17] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[17] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[17].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[17].Id[1]  =  17      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[17].put(sys_operation_lane[17])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[17].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[17];                                                                                                                
            join_none                                                                                                                             
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[18] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[18] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[18].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[18].Id[1]  =  18      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[18].put(sys_operation_lane[18])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[18].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[18];                                                                                                                
            join_none                                                                                                                             
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[19] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[19] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[19].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[19].Id[1]  =  19      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[19].put(sys_operation_lane[19])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[19].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[19];                                                                                                                
            join_none                                                                                                                             
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[20] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[20] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[20].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[20].Id[1]  =  20      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[20].put(sys_operation_lane[20])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[20].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[20];                                                                                                                
            join_none                                                                                                                             
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[21] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[21] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[21].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[21].Id[1]  =  21      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[21].put(sys_operation_lane[21])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[21].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[21];                                                                                                                
            join_none                                                                                                                             
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[22] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[22] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[22].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[22].Id[1]  =  22      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[22].put(sys_operation_lane[22])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[22].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[22];                                                                                                                
            join_none                                                                                                                             
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[23] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[23] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[23].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[23].Id[1]  =  23      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[23].put(sys_operation_lane[23])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[23].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[23];                                                                                                                
            join_none                                                                                                                             
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[24] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[24] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[24].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[24].Id[1]  =  24      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[24].put(sys_operation_lane[24])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[24].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[24];                                                                                                                
            join_none                                                                                                                             
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[25] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[25] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[25].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[25].Id[1]  =  25      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[25].put(sys_operation_lane[25])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[25].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[25];                                                                                                                
            join_none                                                                                                                             
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[26] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[26] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[26].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[26].Id[1]  =  26      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[26].put(sys_operation_lane[26])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[26].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[26];                                                                                                                
            join_none                                                                                                                             
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[27] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[27] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[27].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[27].Id[1]  =  27      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[27].put(sys_operation_lane[27])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[27].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[27];                                                                                                                
            join_none                                                                                                                             
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[28] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[28] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[28].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[28].Id[1]  =  28      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[28].put(sys_operation_lane[28])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[28].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[28];                                                                                                                
            join_none                                                                                                                             
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[29] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[29] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[29].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[29].Id[1]  =  29      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[29].put(sys_operation_lane[29])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[29].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[29];                                                                                                                
            join_none                                                                                                                             
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[30] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[30] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[30].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[30].Id[1]  =  30      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[30].put(sys_operation_lane[30])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[30].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[30];                                                                                                                
            join_none                                                                                                                             
            fork                                                                                                                                  
                // Making sure we create new operand arrays using a deep copy method doesnt seem to be neccessary, but do it anyway (flaky SV)    
                //sys_operation_lane[31] = new sys_operation_mgr ;                                                                               
                // base_operation deep copy also reseeds RNG                                                                                      
                sys_operation_lane[31] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                // The copy copies RNG so need to reseed otherwise we will create the same contents for each lane                                 
                // sys_operation_lane[31].srandom($urandom)       ; // done by deep copy routine                                                 
                sys_operation_lane[31].Id[1]  =  31      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                mgr2gen[31].put(sys_operation_lane[31])                    ;                                                                    
                                                                                                                                                  
                // DEBUG                                                                                                                          
                /*                                                                                                                                
                if (this.Id == 63)                                                                                                                
                  begin                                                                                                                           
                    sys_operation_lane[31].displayOperation();                                                                                   
                  end                                                                                                                             
                */                                                                                                                                
                // now wait for generator                                                                                                         
                @mgr2gen_ack[31];                                                                                                                
            join_none                                                                                                                             
