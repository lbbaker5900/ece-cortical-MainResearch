
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe0__stu__valid        ( UpstreamStackBus[0].pe__stu__valid             ),      
        .pe0__stu__cntl         ( UpstreamStackBus[0].pe__stu__cntl              ),      
        .stu__pe0__ready        ( 1'b1                                            ),      
        //.stu__pe0__ready        ( UpstreamStackBus[0].stu__pe__ready     ),      
        .pe0__stu__type         ( UpstreamStackBus[0].pe__stu__type              ),      
        .pe0__stu__data         ( UpstreamStackBus[0].pe__stu__data              ),      
        .pe0__stu__oob_data     ( UpstreamStackBus[0].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe1__stu__valid        ( UpstreamStackBus[1].pe__stu__valid             ),      
        .pe1__stu__cntl         ( UpstreamStackBus[1].pe__stu__cntl              ),      
        .stu__pe1__ready        ( 1'b1                                            ),      
        //.stu__pe1__ready        ( UpstreamStackBus[1].stu__pe__ready     ),      
        .pe1__stu__type         ( UpstreamStackBus[1].pe__stu__type              ),      
        .pe1__stu__data         ( UpstreamStackBus[1].pe__stu__data              ),      
        .pe1__stu__oob_data     ( UpstreamStackBus[1].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe2__stu__valid        ( UpstreamStackBus[2].pe__stu__valid             ),      
        .pe2__stu__cntl         ( UpstreamStackBus[2].pe__stu__cntl              ),      
        .stu__pe2__ready        ( 1'b1                                            ),      
        //.stu__pe2__ready        ( UpstreamStackBus[2].stu__pe__ready     ),      
        .pe2__stu__type         ( UpstreamStackBus[2].pe__stu__type              ),      
        .pe2__stu__data         ( UpstreamStackBus[2].pe__stu__data              ),      
        .pe2__stu__oob_data     ( UpstreamStackBus[2].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe3__stu__valid        ( UpstreamStackBus[3].pe__stu__valid             ),      
        .pe3__stu__cntl         ( UpstreamStackBus[3].pe__stu__cntl              ),      
        .stu__pe3__ready        ( 1'b1                                            ),      
        //.stu__pe3__ready        ( UpstreamStackBus[3].stu__pe__ready     ),      
        .pe3__stu__type         ( UpstreamStackBus[3].pe__stu__type              ),      
        .pe3__stu__data         ( UpstreamStackBus[3].pe__stu__data              ),      
        .pe3__stu__oob_data     ( UpstreamStackBus[3].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe4__stu__valid        ( UpstreamStackBus[4].pe__stu__valid             ),      
        .pe4__stu__cntl         ( UpstreamStackBus[4].pe__stu__cntl              ),      
        .stu__pe4__ready        ( 1'b1                                            ),      
        //.stu__pe4__ready        ( UpstreamStackBus[4].stu__pe__ready     ),      
        .pe4__stu__type         ( UpstreamStackBus[4].pe__stu__type              ),      
        .pe4__stu__data         ( UpstreamStackBus[4].pe__stu__data              ),      
        .pe4__stu__oob_data     ( UpstreamStackBus[4].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe5__stu__valid        ( UpstreamStackBus[5].pe__stu__valid             ),      
        .pe5__stu__cntl         ( UpstreamStackBus[5].pe__stu__cntl              ),      
        .stu__pe5__ready        ( 1'b1                                            ),      
        //.stu__pe5__ready        ( UpstreamStackBus[5].stu__pe__ready     ),      
        .pe5__stu__type         ( UpstreamStackBus[5].pe__stu__type              ),      
        .pe5__stu__data         ( UpstreamStackBus[5].pe__stu__data              ),      
        .pe5__stu__oob_data     ( UpstreamStackBus[5].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe6__stu__valid        ( UpstreamStackBus[6].pe__stu__valid             ),      
        .pe6__stu__cntl         ( UpstreamStackBus[6].pe__stu__cntl              ),      
        .stu__pe6__ready        ( 1'b1                                            ),      
        //.stu__pe6__ready        ( UpstreamStackBus[6].stu__pe__ready     ),      
        .pe6__stu__type         ( UpstreamStackBus[6].pe__stu__type              ),      
        .pe6__stu__data         ( UpstreamStackBus[6].pe__stu__data              ),      
        .pe6__stu__oob_data     ( UpstreamStackBus[6].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe7__stu__valid        ( UpstreamStackBus[7].pe__stu__valid             ),      
        .pe7__stu__cntl         ( UpstreamStackBus[7].pe__stu__cntl              ),      
        .stu__pe7__ready        ( 1'b1                                            ),      
        //.stu__pe7__ready        ( UpstreamStackBus[7].stu__pe__ready     ),      
        .pe7__stu__type         ( UpstreamStackBus[7].pe__stu__type              ),      
        .pe7__stu__data         ( UpstreamStackBus[7].pe__stu__data              ),      
        .pe7__stu__oob_data     ( UpstreamStackBus[7].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe8__stu__valid        ( UpstreamStackBus[8].pe__stu__valid             ),      
        .pe8__stu__cntl         ( UpstreamStackBus[8].pe__stu__cntl              ),      
        .stu__pe8__ready        ( 1'b1                                            ),      
        //.stu__pe8__ready        ( UpstreamStackBus[8].stu__pe__ready     ),      
        .pe8__stu__type         ( UpstreamStackBus[8].pe__stu__type              ),      
        .pe8__stu__data         ( UpstreamStackBus[8].pe__stu__data              ),      
        .pe8__stu__oob_data     ( UpstreamStackBus[8].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe9__stu__valid        ( UpstreamStackBus[9].pe__stu__valid             ),      
        .pe9__stu__cntl         ( UpstreamStackBus[9].pe__stu__cntl              ),      
        .stu__pe9__ready        ( 1'b1                                            ),      
        //.stu__pe9__ready        ( UpstreamStackBus[9].stu__pe__ready     ),      
        .pe9__stu__type         ( UpstreamStackBus[9].pe__stu__type              ),      
        .pe9__stu__data         ( UpstreamStackBus[9].pe__stu__data              ),      
        .pe9__stu__oob_data     ( UpstreamStackBus[9].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe10__stu__valid        ( UpstreamStackBus[10].pe__stu__valid             ),      
        .pe10__stu__cntl         ( UpstreamStackBus[10].pe__stu__cntl              ),      
        .stu__pe10__ready        ( 1'b1                                            ),      
        //.stu__pe10__ready        ( UpstreamStackBus[10].stu__pe__ready     ),      
        .pe10__stu__type         ( UpstreamStackBus[10].pe__stu__type              ),      
        .pe10__stu__data         ( UpstreamStackBus[10].pe__stu__data              ),      
        .pe10__stu__oob_data     ( UpstreamStackBus[10].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe11__stu__valid        ( UpstreamStackBus[11].pe__stu__valid             ),      
        .pe11__stu__cntl         ( UpstreamStackBus[11].pe__stu__cntl              ),      
        .stu__pe11__ready        ( 1'b1                                            ),      
        //.stu__pe11__ready        ( UpstreamStackBus[11].stu__pe__ready     ),      
        .pe11__stu__type         ( UpstreamStackBus[11].pe__stu__type              ),      
        .pe11__stu__data         ( UpstreamStackBus[11].pe__stu__data              ),      
        .pe11__stu__oob_data     ( UpstreamStackBus[11].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe12__stu__valid        ( UpstreamStackBus[12].pe__stu__valid             ),      
        .pe12__stu__cntl         ( UpstreamStackBus[12].pe__stu__cntl              ),      
        .stu__pe12__ready        ( 1'b1                                            ),      
        //.stu__pe12__ready        ( UpstreamStackBus[12].stu__pe__ready     ),      
        .pe12__stu__type         ( UpstreamStackBus[12].pe__stu__type              ),      
        .pe12__stu__data         ( UpstreamStackBus[12].pe__stu__data              ),      
        .pe12__stu__oob_data     ( UpstreamStackBus[12].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe13__stu__valid        ( UpstreamStackBus[13].pe__stu__valid             ),      
        .pe13__stu__cntl         ( UpstreamStackBus[13].pe__stu__cntl              ),      
        .stu__pe13__ready        ( 1'b1                                            ),      
        //.stu__pe13__ready        ( UpstreamStackBus[13].stu__pe__ready     ),      
        .pe13__stu__type         ( UpstreamStackBus[13].pe__stu__type              ),      
        .pe13__stu__data         ( UpstreamStackBus[13].pe__stu__data              ),      
        .pe13__stu__oob_data     ( UpstreamStackBus[13].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe14__stu__valid        ( UpstreamStackBus[14].pe__stu__valid             ),      
        .pe14__stu__cntl         ( UpstreamStackBus[14].pe__stu__cntl              ),      
        .stu__pe14__ready        ( 1'b1                                            ),      
        //.stu__pe14__ready        ( UpstreamStackBus[14].stu__pe__ready     ),      
        .pe14__stu__type         ( UpstreamStackBus[14].pe__stu__type              ),      
        .pe14__stu__data         ( UpstreamStackBus[14].pe__stu__data              ),      
        .pe14__stu__oob_data     ( UpstreamStackBus[14].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe15__stu__valid        ( UpstreamStackBus[15].pe__stu__valid             ),      
        .pe15__stu__cntl         ( UpstreamStackBus[15].pe__stu__cntl              ),      
        .stu__pe15__ready        ( 1'b1                                            ),      
        //.stu__pe15__ready        ( UpstreamStackBus[15].stu__pe__ready     ),      
        .pe15__stu__type         ( UpstreamStackBus[15].pe__stu__type              ),      
        .pe15__stu__data         ( UpstreamStackBus[15].pe__stu__data              ),      
        .pe15__stu__oob_data     ( UpstreamStackBus[15].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe16__stu__valid        ( UpstreamStackBus[16].pe__stu__valid             ),      
        .pe16__stu__cntl         ( UpstreamStackBus[16].pe__stu__cntl              ),      
        .stu__pe16__ready        ( 1'b1                                            ),      
        //.stu__pe16__ready        ( UpstreamStackBus[16].stu__pe__ready     ),      
        .pe16__stu__type         ( UpstreamStackBus[16].pe__stu__type              ),      
        .pe16__stu__data         ( UpstreamStackBus[16].pe__stu__data              ),      
        .pe16__stu__oob_data     ( UpstreamStackBus[16].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe17__stu__valid        ( UpstreamStackBus[17].pe__stu__valid             ),      
        .pe17__stu__cntl         ( UpstreamStackBus[17].pe__stu__cntl              ),      
        .stu__pe17__ready        ( 1'b1                                            ),      
        //.stu__pe17__ready        ( UpstreamStackBus[17].stu__pe__ready     ),      
        .pe17__stu__type         ( UpstreamStackBus[17].pe__stu__type              ),      
        .pe17__stu__data         ( UpstreamStackBus[17].pe__stu__data              ),      
        .pe17__stu__oob_data     ( UpstreamStackBus[17].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe18__stu__valid        ( UpstreamStackBus[18].pe__stu__valid             ),      
        .pe18__stu__cntl         ( UpstreamStackBus[18].pe__stu__cntl              ),      
        .stu__pe18__ready        ( 1'b1                                            ),      
        //.stu__pe18__ready        ( UpstreamStackBus[18].stu__pe__ready     ),      
        .pe18__stu__type         ( UpstreamStackBus[18].pe__stu__type              ),      
        .pe18__stu__data         ( UpstreamStackBus[18].pe__stu__data              ),      
        .pe18__stu__oob_data     ( UpstreamStackBus[18].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe19__stu__valid        ( UpstreamStackBus[19].pe__stu__valid             ),      
        .pe19__stu__cntl         ( UpstreamStackBus[19].pe__stu__cntl              ),      
        .stu__pe19__ready        ( 1'b1                                            ),      
        //.stu__pe19__ready        ( UpstreamStackBus[19].stu__pe__ready     ),      
        .pe19__stu__type         ( UpstreamStackBus[19].pe__stu__type              ),      
        .pe19__stu__data         ( UpstreamStackBus[19].pe__stu__data              ),      
        .pe19__stu__oob_data     ( UpstreamStackBus[19].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe20__stu__valid        ( UpstreamStackBus[20].pe__stu__valid             ),      
        .pe20__stu__cntl         ( UpstreamStackBus[20].pe__stu__cntl              ),      
        .stu__pe20__ready        ( 1'b1                                            ),      
        //.stu__pe20__ready        ( UpstreamStackBus[20].stu__pe__ready     ),      
        .pe20__stu__type         ( UpstreamStackBus[20].pe__stu__type              ),      
        .pe20__stu__data         ( UpstreamStackBus[20].pe__stu__data              ),      
        .pe20__stu__oob_data     ( UpstreamStackBus[20].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe21__stu__valid        ( UpstreamStackBus[21].pe__stu__valid             ),      
        .pe21__stu__cntl         ( UpstreamStackBus[21].pe__stu__cntl              ),      
        .stu__pe21__ready        ( 1'b1                                            ),      
        //.stu__pe21__ready        ( UpstreamStackBus[21].stu__pe__ready     ),      
        .pe21__stu__type         ( UpstreamStackBus[21].pe__stu__type              ),      
        .pe21__stu__data         ( UpstreamStackBus[21].pe__stu__data              ),      
        .pe21__stu__oob_data     ( UpstreamStackBus[21].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe22__stu__valid        ( UpstreamStackBus[22].pe__stu__valid             ),      
        .pe22__stu__cntl         ( UpstreamStackBus[22].pe__stu__cntl              ),      
        .stu__pe22__ready        ( 1'b1                                            ),      
        //.stu__pe22__ready        ( UpstreamStackBus[22].stu__pe__ready     ),      
        .pe22__stu__type         ( UpstreamStackBus[22].pe__stu__type              ),      
        .pe22__stu__data         ( UpstreamStackBus[22].pe__stu__data              ),      
        .pe22__stu__oob_data     ( UpstreamStackBus[22].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe23__stu__valid        ( UpstreamStackBus[23].pe__stu__valid             ),      
        .pe23__stu__cntl         ( UpstreamStackBus[23].pe__stu__cntl              ),      
        .stu__pe23__ready        ( 1'b1                                            ),      
        //.stu__pe23__ready        ( UpstreamStackBus[23].stu__pe__ready     ),      
        .pe23__stu__type         ( UpstreamStackBus[23].pe__stu__type              ),      
        .pe23__stu__data         ( UpstreamStackBus[23].pe__stu__data              ),      
        .pe23__stu__oob_data     ( UpstreamStackBus[23].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe24__stu__valid        ( UpstreamStackBus[24].pe__stu__valid             ),      
        .pe24__stu__cntl         ( UpstreamStackBus[24].pe__stu__cntl              ),      
        .stu__pe24__ready        ( 1'b1                                            ),      
        //.stu__pe24__ready        ( UpstreamStackBus[24].stu__pe__ready     ),      
        .pe24__stu__type         ( UpstreamStackBus[24].pe__stu__type              ),      
        .pe24__stu__data         ( UpstreamStackBus[24].pe__stu__data              ),      
        .pe24__stu__oob_data     ( UpstreamStackBus[24].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe25__stu__valid        ( UpstreamStackBus[25].pe__stu__valid             ),      
        .pe25__stu__cntl         ( UpstreamStackBus[25].pe__stu__cntl              ),      
        .stu__pe25__ready        ( 1'b1                                            ),      
        //.stu__pe25__ready        ( UpstreamStackBus[25].stu__pe__ready     ),      
        .pe25__stu__type         ( UpstreamStackBus[25].pe__stu__type              ),      
        .pe25__stu__data         ( UpstreamStackBus[25].pe__stu__data              ),      
        .pe25__stu__oob_data     ( UpstreamStackBus[25].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe26__stu__valid        ( UpstreamStackBus[26].pe__stu__valid             ),      
        .pe26__stu__cntl         ( UpstreamStackBus[26].pe__stu__cntl              ),      
        .stu__pe26__ready        ( 1'b1                                            ),      
        //.stu__pe26__ready        ( UpstreamStackBus[26].stu__pe__ready     ),      
        .pe26__stu__type         ( UpstreamStackBus[26].pe__stu__type              ),      
        .pe26__stu__data         ( UpstreamStackBus[26].pe__stu__data              ),      
        .pe26__stu__oob_data     ( UpstreamStackBus[26].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe27__stu__valid        ( UpstreamStackBus[27].pe__stu__valid             ),      
        .pe27__stu__cntl         ( UpstreamStackBus[27].pe__stu__cntl              ),      
        .stu__pe27__ready        ( 1'b1                                            ),      
        //.stu__pe27__ready        ( UpstreamStackBus[27].stu__pe__ready     ),      
        .pe27__stu__type         ( UpstreamStackBus[27].pe__stu__type              ),      
        .pe27__stu__data         ( UpstreamStackBus[27].pe__stu__data              ),      
        .pe27__stu__oob_data     ( UpstreamStackBus[27].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe28__stu__valid        ( UpstreamStackBus[28].pe__stu__valid             ),      
        .pe28__stu__cntl         ( UpstreamStackBus[28].pe__stu__cntl              ),      
        .stu__pe28__ready        ( 1'b1                                            ),      
        //.stu__pe28__ready        ( UpstreamStackBus[28].stu__pe__ready     ),      
        .pe28__stu__type         ( UpstreamStackBus[28].pe__stu__type              ),      
        .pe28__stu__data         ( UpstreamStackBus[28].pe__stu__data              ),      
        .pe28__stu__oob_data     ( UpstreamStackBus[28].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe29__stu__valid        ( UpstreamStackBus[29].pe__stu__valid             ),      
        .pe29__stu__cntl         ( UpstreamStackBus[29].pe__stu__cntl              ),      
        .stu__pe29__ready        ( 1'b1                                            ),      
        //.stu__pe29__ready        ( UpstreamStackBus[29].stu__pe__ready     ),      
        .pe29__stu__type         ( UpstreamStackBus[29].pe__stu__type              ),      
        .pe29__stu__data         ( UpstreamStackBus[29].pe__stu__data              ),      
        .pe29__stu__oob_data     ( UpstreamStackBus[29].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe30__stu__valid        ( UpstreamStackBus[30].pe__stu__valid             ),      
        .pe30__stu__cntl         ( UpstreamStackBus[30].pe__stu__cntl              ),      
        .stu__pe30__ready        ( 1'b1                                            ),      
        //.stu__pe30__ready        ( UpstreamStackBus[30].stu__pe__ready     ),      
        .pe30__stu__type         ( UpstreamStackBus[30].pe__stu__type              ),      
        .pe30__stu__data         ( UpstreamStackBus[30].pe__stu__data              ),      
        .pe30__stu__oob_data     ( UpstreamStackBus[30].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe31__stu__valid        ( UpstreamStackBus[31].pe__stu__valid             ),      
        .pe31__stu__cntl         ( UpstreamStackBus[31].pe__stu__cntl              ),      
        .stu__pe31__ready        ( 1'b1                                            ),      
        //.stu__pe31__ready        ( UpstreamStackBus[31].stu__pe__ready     ),      
        .pe31__stu__type         ( UpstreamStackBus[31].pe__stu__type              ),      
        .pe31__stu__data         ( UpstreamStackBus[31].pe__stu__data              ),      
        .pe31__stu__oob_data     ( UpstreamStackBus[31].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe32__stu__valid        ( UpstreamStackBus[32].pe__stu__valid             ),      
        .pe32__stu__cntl         ( UpstreamStackBus[32].pe__stu__cntl              ),      
        .stu__pe32__ready        ( 1'b1                                            ),      
        //.stu__pe32__ready        ( UpstreamStackBus[32].stu__pe__ready     ),      
        .pe32__stu__type         ( UpstreamStackBus[32].pe__stu__type              ),      
        .pe32__stu__data         ( UpstreamStackBus[32].pe__stu__data              ),      
        .pe32__stu__oob_data     ( UpstreamStackBus[32].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe33__stu__valid        ( UpstreamStackBus[33].pe__stu__valid             ),      
        .pe33__stu__cntl         ( UpstreamStackBus[33].pe__stu__cntl              ),      
        .stu__pe33__ready        ( 1'b1                                            ),      
        //.stu__pe33__ready        ( UpstreamStackBus[33].stu__pe__ready     ),      
        .pe33__stu__type         ( UpstreamStackBus[33].pe__stu__type              ),      
        .pe33__stu__data         ( UpstreamStackBus[33].pe__stu__data              ),      
        .pe33__stu__oob_data     ( UpstreamStackBus[33].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe34__stu__valid        ( UpstreamStackBus[34].pe__stu__valid             ),      
        .pe34__stu__cntl         ( UpstreamStackBus[34].pe__stu__cntl              ),      
        .stu__pe34__ready        ( 1'b1                                            ),      
        //.stu__pe34__ready        ( UpstreamStackBus[34].stu__pe__ready     ),      
        .pe34__stu__type         ( UpstreamStackBus[34].pe__stu__type              ),      
        .pe34__stu__data         ( UpstreamStackBus[34].pe__stu__data              ),      
        .pe34__stu__oob_data     ( UpstreamStackBus[34].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe35__stu__valid        ( UpstreamStackBus[35].pe__stu__valid             ),      
        .pe35__stu__cntl         ( UpstreamStackBus[35].pe__stu__cntl              ),      
        .stu__pe35__ready        ( 1'b1                                            ),      
        //.stu__pe35__ready        ( UpstreamStackBus[35].stu__pe__ready     ),      
        .pe35__stu__type         ( UpstreamStackBus[35].pe__stu__type              ),      
        .pe35__stu__data         ( UpstreamStackBus[35].pe__stu__data              ),      
        .pe35__stu__oob_data     ( UpstreamStackBus[35].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe36__stu__valid        ( UpstreamStackBus[36].pe__stu__valid             ),      
        .pe36__stu__cntl         ( UpstreamStackBus[36].pe__stu__cntl              ),      
        .stu__pe36__ready        ( 1'b1                                            ),      
        //.stu__pe36__ready        ( UpstreamStackBus[36].stu__pe__ready     ),      
        .pe36__stu__type         ( UpstreamStackBus[36].pe__stu__type              ),      
        .pe36__stu__data         ( UpstreamStackBus[36].pe__stu__data              ),      
        .pe36__stu__oob_data     ( UpstreamStackBus[36].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe37__stu__valid        ( UpstreamStackBus[37].pe__stu__valid             ),      
        .pe37__stu__cntl         ( UpstreamStackBus[37].pe__stu__cntl              ),      
        .stu__pe37__ready        ( 1'b1                                            ),      
        //.stu__pe37__ready        ( UpstreamStackBus[37].stu__pe__ready     ),      
        .pe37__stu__type         ( UpstreamStackBus[37].pe__stu__type              ),      
        .pe37__stu__data         ( UpstreamStackBus[37].pe__stu__data              ),      
        .pe37__stu__oob_data     ( UpstreamStackBus[37].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe38__stu__valid        ( UpstreamStackBus[38].pe__stu__valid             ),      
        .pe38__stu__cntl         ( UpstreamStackBus[38].pe__stu__cntl              ),      
        .stu__pe38__ready        ( 1'b1                                            ),      
        //.stu__pe38__ready        ( UpstreamStackBus[38].stu__pe__ready     ),      
        .pe38__stu__type         ( UpstreamStackBus[38].pe__stu__type              ),      
        .pe38__stu__data         ( UpstreamStackBus[38].pe__stu__data              ),      
        .pe38__stu__oob_data     ( UpstreamStackBus[38].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe39__stu__valid        ( UpstreamStackBus[39].pe__stu__valid             ),      
        .pe39__stu__cntl         ( UpstreamStackBus[39].pe__stu__cntl              ),      
        .stu__pe39__ready        ( 1'b1                                            ),      
        //.stu__pe39__ready        ( UpstreamStackBus[39].stu__pe__ready     ),      
        .pe39__stu__type         ( UpstreamStackBus[39].pe__stu__type              ),      
        .pe39__stu__data         ( UpstreamStackBus[39].pe__stu__data              ),      
        .pe39__stu__oob_data     ( UpstreamStackBus[39].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe40__stu__valid        ( UpstreamStackBus[40].pe__stu__valid             ),      
        .pe40__stu__cntl         ( UpstreamStackBus[40].pe__stu__cntl              ),      
        .stu__pe40__ready        ( 1'b1                                            ),      
        //.stu__pe40__ready        ( UpstreamStackBus[40].stu__pe__ready     ),      
        .pe40__stu__type         ( UpstreamStackBus[40].pe__stu__type              ),      
        .pe40__stu__data         ( UpstreamStackBus[40].pe__stu__data              ),      
        .pe40__stu__oob_data     ( UpstreamStackBus[40].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe41__stu__valid        ( UpstreamStackBus[41].pe__stu__valid             ),      
        .pe41__stu__cntl         ( UpstreamStackBus[41].pe__stu__cntl              ),      
        .stu__pe41__ready        ( 1'b1                                            ),      
        //.stu__pe41__ready        ( UpstreamStackBus[41].stu__pe__ready     ),      
        .pe41__stu__type         ( UpstreamStackBus[41].pe__stu__type              ),      
        .pe41__stu__data         ( UpstreamStackBus[41].pe__stu__data              ),      
        .pe41__stu__oob_data     ( UpstreamStackBus[41].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe42__stu__valid        ( UpstreamStackBus[42].pe__stu__valid             ),      
        .pe42__stu__cntl         ( UpstreamStackBus[42].pe__stu__cntl              ),      
        .stu__pe42__ready        ( 1'b1                                            ),      
        //.stu__pe42__ready        ( UpstreamStackBus[42].stu__pe__ready     ),      
        .pe42__stu__type         ( UpstreamStackBus[42].pe__stu__type              ),      
        .pe42__stu__data         ( UpstreamStackBus[42].pe__stu__data              ),      
        .pe42__stu__oob_data     ( UpstreamStackBus[42].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe43__stu__valid        ( UpstreamStackBus[43].pe__stu__valid             ),      
        .pe43__stu__cntl         ( UpstreamStackBus[43].pe__stu__cntl              ),      
        .stu__pe43__ready        ( 1'b1                                            ),      
        //.stu__pe43__ready        ( UpstreamStackBus[43].stu__pe__ready     ),      
        .pe43__stu__type         ( UpstreamStackBus[43].pe__stu__type              ),      
        .pe43__stu__data         ( UpstreamStackBus[43].pe__stu__data              ),      
        .pe43__stu__oob_data     ( UpstreamStackBus[43].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe44__stu__valid        ( UpstreamStackBus[44].pe__stu__valid             ),      
        .pe44__stu__cntl         ( UpstreamStackBus[44].pe__stu__cntl              ),      
        .stu__pe44__ready        ( 1'b1                                            ),      
        //.stu__pe44__ready        ( UpstreamStackBus[44].stu__pe__ready     ),      
        .pe44__stu__type         ( UpstreamStackBus[44].pe__stu__type              ),      
        .pe44__stu__data         ( UpstreamStackBus[44].pe__stu__data              ),      
        .pe44__stu__oob_data     ( UpstreamStackBus[44].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe45__stu__valid        ( UpstreamStackBus[45].pe__stu__valid             ),      
        .pe45__stu__cntl         ( UpstreamStackBus[45].pe__stu__cntl              ),      
        .stu__pe45__ready        ( 1'b1                                            ),      
        //.stu__pe45__ready        ( UpstreamStackBus[45].stu__pe__ready     ),      
        .pe45__stu__type         ( UpstreamStackBus[45].pe__stu__type              ),      
        .pe45__stu__data         ( UpstreamStackBus[45].pe__stu__data              ),      
        .pe45__stu__oob_data     ( UpstreamStackBus[45].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe46__stu__valid        ( UpstreamStackBus[46].pe__stu__valid             ),      
        .pe46__stu__cntl         ( UpstreamStackBus[46].pe__stu__cntl              ),      
        .stu__pe46__ready        ( 1'b1                                            ),      
        //.stu__pe46__ready        ( UpstreamStackBus[46].stu__pe__ready     ),      
        .pe46__stu__type         ( UpstreamStackBus[46].pe__stu__type              ),      
        .pe46__stu__data         ( UpstreamStackBus[46].pe__stu__data              ),      
        .pe46__stu__oob_data     ( UpstreamStackBus[46].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe47__stu__valid        ( UpstreamStackBus[47].pe__stu__valid             ),      
        .pe47__stu__cntl         ( UpstreamStackBus[47].pe__stu__cntl              ),      
        .stu__pe47__ready        ( 1'b1                                            ),      
        //.stu__pe47__ready        ( UpstreamStackBus[47].stu__pe__ready     ),      
        .pe47__stu__type         ( UpstreamStackBus[47].pe__stu__type              ),      
        .pe47__stu__data         ( UpstreamStackBus[47].pe__stu__data              ),      
        .pe47__stu__oob_data     ( UpstreamStackBus[47].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe48__stu__valid        ( UpstreamStackBus[48].pe__stu__valid             ),      
        .pe48__stu__cntl         ( UpstreamStackBus[48].pe__stu__cntl              ),      
        .stu__pe48__ready        ( 1'b1                                            ),      
        //.stu__pe48__ready        ( UpstreamStackBus[48].stu__pe__ready     ),      
        .pe48__stu__type         ( UpstreamStackBus[48].pe__stu__type              ),      
        .pe48__stu__data         ( UpstreamStackBus[48].pe__stu__data              ),      
        .pe48__stu__oob_data     ( UpstreamStackBus[48].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe49__stu__valid        ( UpstreamStackBus[49].pe__stu__valid             ),      
        .pe49__stu__cntl         ( UpstreamStackBus[49].pe__stu__cntl              ),      
        .stu__pe49__ready        ( 1'b1                                            ),      
        //.stu__pe49__ready        ( UpstreamStackBus[49].stu__pe__ready     ),      
        .pe49__stu__type         ( UpstreamStackBus[49].pe__stu__type              ),      
        .pe49__stu__data         ( UpstreamStackBus[49].pe__stu__data              ),      
        .pe49__stu__oob_data     ( UpstreamStackBus[49].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe50__stu__valid        ( UpstreamStackBus[50].pe__stu__valid             ),      
        .pe50__stu__cntl         ( UpstreamStackBus[50].pe__stu__cntl              ),      
        .stu__pe50__ready        ( 1'b1                                            ),      
        //.stu__pe50__ready        ( UpstreamStackBus[50].stu__pe__ready     ),      
        .pe50__stu__type         ( UpstreamStackBus[50].pe__stu__type              ),      
        .pe50__stu__data         ( UpstreamStackBus[50].pe__stu__data              ),      
        .pe50__stu__oob_data     ( UpstreamStackBus[50].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe51__stu__valid        ( UpstreamStackBus[51].pe__stu__valid             ),      
        .pe51__stu__cntl         ( UpstreamStackBus[51].pe__stu__cntl              ),      
        .stu__pe51__ready        ( 1'b1                                            ),      
        //.stu__pe51__ready        ( UpstreamStackBus[51].stu__pe__ready     ),      
        .pe51__stu__type         ( UpstreamStackBus[51].pe__stu__type              ),      
        .pe51__stu__data         ( UpstreamStackBus[51].pe__stu__data              ),      
        .pe51__stu__oob_data     ( UpstreamStackBus[51].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe52__stu__valid        ( UpstreamStackBus[52].pe__stu__valid             ),      
        .pe52__stu__cntl         ( UpstreamStackBus[52].pe__stu__cntl              ),      
        .stu__pe52__ready        ( 1'b1                                            ),      
        //.stu__pe52__ready        ( UpstreamStackBus[52].stu__pe__ready     ),      
        .pe52__stu__type         ( UpstreamStackBus[52].pe__stu__type              ),      
        .pe52__stu__data         ( UpstreamStackBus[52].pe__stu__data              ),      
        .pe52__stu__oob_data     ( UpstreamStackBus[52].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe53__stu__valid        ( UpstreamStackBus[53].pe__stu__valid             ),      
        .pe53__stu__cntl         ( UpstreamStackBus[53].pe__stu__cntl              ),      
        .stu__pe53__ready        ( 1'b1                                            ),      
        //.stu__pe53__ready        ( UpstreamStackBus[53].stu__pe__ready     ),      
        .pe53__stu__type         ( UpstreamStackBus[53].pe__stu__type              ),      
        .pe53__stu__data         ( UpstreamStackBus[53].pe__stu__data              ),      
        .pe53__stu__oob_data     ( UpstreamStackBus[53].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe54__stu__valid        ( UpstreamStackBus[54].pe__stu__valid             ),      
        .pe54__stu__cntl         ( UpstreamStackBus[54].pe__stu__cntl              ),      
        .stu__pe54__ready        ( 1'b1                                            ),      
        //.stu__pe54__ready        ( UpstreamStackBus[54].stu__pe__ready     ),      
        .pe54__stu__type         ( UpstreamStackBus[54].pe__stu__type              ),      
        .pe54__stu__data         ( UpstreamStackBus[54].pe__stu__data              ),      
        .pe54__stu__oob_data     ( UpstreamStackBus[54].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe55__stu__valid        ( UpstreamStackBus[55].pe__stu__valid             ),      
        .pe55__stu__cntl         ( UpstreamStackBus[55].pe__stu__cntl              ),      
        .stu__pe55__ready        ( 1'b1                                            ),      
        //.stu__pe55__ready        ( UpstreamStackBus[55].stu__pe__ready     ),      
        .pe55__stu__type         ( UpstreamStackBus[55].pe__stu__type              ),      
        .pe55__stu__data         ( UpstreamStackBus[55].pe__stu__data              ),      
        .pe55__stu__oob_data     ( UpstreamStackBus[55].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe56__stu__valid        ( UpstreamStackBus[56].pe__stu__valid             ),      
        .pe56__stu__cntl         ( UpstreamStackBus[56].pe__stu__cntl              ),      
        .stu__pe56__ready        ( 1'b1                                            ),      
        //.stu__pe56__ready        ( UpstreamStackBus[56].stu__pe__ready     ),      
        .pe56__stu__type         ( UpstreamStackBus[56].pe__stu__type              ),      
        .pe56__stu__data         ( UpstreamStackBus[56].pe__stu__data              ),      
        .pe56__stu__oob_data     ( UpstreamStackBus[56].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe57__stu__valid        ( UpstreamStackBus[57].pe__stu__valid             ),      
        .pe57__stu__cntl         ( UpstreamStackBus[57].pe__stu__cntl              ),      
        .stu__pe57__ready        ( 1'b1                                            ),      
        //.stu__pe57__ready        ( UpstreamStackBus[57].stu__pe__ready     ),      
        .pe57__stu__type         ( UpstreamStackBus[57].pe__stu__type              ),      
        .pe57__stu__data         ( UpstreamStackBus[57].pe__stu__data              ),      
        .pe57__stu__oob_data     ( UpstreamStackBus[57].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe58__stu__valid        ( UpstreamStackBus[58].pe__stu__valid             ),      
        .pe58__stu__cntl         ( UpstreamStackBus[58].pe__stu__cntl              ),      
        .stu__pe58__ready        ( 1'b1                                            ),      
        //.stu__pe58__ready        ( UpstreamStackBus[58].stu__pe__ready     ),      
        .pe58__stu__type         ( UpstreamStackBus[58].pe__stu__type              ),      
        .pe58__stu__data         ( UpstreamStackBus[58].pe__stu__data              ),      
        .pe58__stu__oob_data     ( UpstreamStackBus[58].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe59__stu__valid        ( UpstreamStackBus[59].pe__stu__valid             ),      
        .pe59__stu__cntl         ( UpstreamStackBus[59].pe__stu__cntl              ),      
        .stu__pe59__ready        ( 1'b1                                            ),      
        //.stu__pe59__ready        ( UpstreamStackBus[59].stu__pe__ready     ),      
        .pe59__stu__type         ( UpstreamStackBus[59].pe__stu__type              ),      
        .pe59__stu__data         ( UpstreamStackBus[59].pe__stu__data              ),      
        .pe59__stu__oob_data     ( UpstreamStackBus[59].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe60__stu__valid        ( UpstreamStackBus[60].pe__stu__valid             ),      
        .pe60__stu__cntl         ( UpstreamStackBus[60].pe__stu__cntl              ),      
        .stu__pe60__ready        ( 1'b1                                            ),      
        //.stu__pe60__ready        ( UpstreamStackBus[60].stu__pe__ready     ),      
        .pe60__stu__type         ( UpstreamStackBus[60].pe__stu__type              ),      
        .pe60__stu__data         ( UpstreamStackBus[60].pe__stu__data              ),      
        .pe60__stu__oob_data     ( UpstreamStackBus[60].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe61__stu__valid        ( UpstreamStackBus[61].pe__stu__valid             ),      
        .pe61__stu__cntl         ( UpstreamStackBus[61].pe__stu__cntl              ),      
        .stu__pe61__ready        ( 1'b1                                            ),      
        //.stu__pe61__ready        ( UpstreamStackBus[61].stu__pe__ready     ),      
        .pe61__stu__type         ( UpstreamStackBus[61].pe__stu__type              ),      
        .pe61__stu__data         ( UpstreamStackBus[61].pe__stu__data              ),      
        .pe61__stu__oob_data     ( UpstreamStackBus[61].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe62__stu__valid        ( UpstreamStackBus[62].pe__stu__valid             ),      
        .pe62__stu__cntl         ( UpstreamStackBus[62].pe__stu__cntl              ),      
        .stu__pe62__ready        ( 1'b1                                            ),      
        //.stu__pe62__ready        ( UpstreamStackBus[62].stu__pe__ready     ),      
        .pe62__stu__type         ( UpstreamStackBus[62].pe__stu__type              ),      
        .pe62__stu__data         ( UpstreamStackBus[62].pe__stu__data              ),      
        .pe62__stu__oob_data     ( UpstreamStackBus[62].pe__stu__oob_data          ),      
        
        //  - doesnt seem to work if you use cb_test for observed signals                                                       
        .pe63__stu__valid        ( UpstreamStackBus[63].pe__stu__valid             ),      
        .pe63__stu__cntl         ( UpstreamStackBus[63].pe__stu__cntl              ),      
        .stu__pe63__ready        ( 1'b1                                            ),      
        //.stu__pe63__ready        ( UpstreamStackBus[63].stu__pe__ready     ),      
        .pe63__stu__type         ( UpstreamStackBus[63].pe__stu__type              ),      
        .pe63__stu__data         ( UpstreamStackBus[63].pe__stu__data              ),      
        .pe63__stu__oob_data     ( UpstreamStackBus[63].pe__stu__oob_data          ),      
        