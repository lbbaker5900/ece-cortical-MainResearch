
//            begin
//              ldst_driver[0].reset()  ;
//            end
//            begin
//              mgr[0].reset()  ;
//            end
//            begin
//              oob_drv[0].reset()  ;
//            end
//            begin
//              up_check[0].reset()  ;
//            end
//            begin
//              gen[0][0].reset()  ;
//            end
//            begin
//              drv[0][0].reset()  ;
//            end
//            begin
//              mem_check[0][0].reset()  ;
//            end
            begin
              rf_driver[0][0].reset()  ;
            end

//            begin
//              gen[0][1].reset()  ;
//            end
//            begin
//              drv[0][1].reset()  ;
//            end
//            begin
//              mem_check[0][1].reset()  ;
//            end
            begin
              rf_driver[0][1].reset()  ;
            end

//            begin
//              gen[0][2].reset()  ;
//            end
//            begin
//              drv[0][2].reset()  ;
//            end
//            begin
//              mem_check[0][2].reset()  ;
//            end
            begin
              rf_driver[0][2].reset()  ;
            end

//            begin
//              gen[0][3].reset()  ;
//            end
//            begin
//              drv[0][3].reset()  ;
//            end
//            begin
//              mem_check[0][3].reset()  ;
//            end
            begin
              rf_driver[0][3].reset()  ;
            end

//            begin
//              gen[0][4].reset()  ;
//            end
//            begin
//              drv[0][4].reset()  ;
//            end
//            begin
//              mem_check[0][4].reset()  ;
//            end
            begin
              rf_driver[0][4].reset()  ;
            end

//            begin
//              gen[0][5].reset()  ;
//            end
//            begin
//              drv[0][5].reset()  ;
//            end
//            begin
//              mem_check[0][5].reset()  ;
//            end
            begin
              rf_driver[0][5].reset()  ;
            end

//            begin
//              gen[0][6].reset()  ;
//            end
//            begin
//              drv[0][6].reset()  ;
//            end
//            begin
//              mem_check[0][6].reset()  ;
//            end
            begin
              rf_driver[0][6].reset()  ;
            end

//            begin
//              gen[0][7].reset()  ;
//            end
//            begin
//              drv[0][7].reset()  ;
//            end
//            begin
//              mem_check[0][7].reset()  ;
//            end
            begin
              rf_driver[0][7].reset()  ;
            end

//            begin
//              gen[0][8].reset()  ;
//            end
//            begin
//              drv[0][8].reset()  ;
//            end
//            begin
//              mem_check[0][8].reset()  ;
//            end
            begin
              rf_driver[0][8].reset()  ;
            end

//            begin
//              gen[0][9].reset()  ;
//            end
//            begin
//              drv[0][9].reset()  ;
//            end
//            begin
//              mem_check[0][9].reset()  ;
//            end
            begin
              rf_driver[0][9].reset()  ;
            end

//            begin
//              gen[0][10].reset()  ;
//            end
//            begin
//              drv[0][10].reset()  ;
//            end
//            begin
//              mem_check[0][10].reset()  ;
//            end
            begin
              rf_driver[0][10].reset()  ;
            end

//            begin
//              gen[0][11].reset()  ;
//            end
//            begin
//              drv[0][11].reset()  ;
//            end
//            begin
//              mem_check[0][11].reset()  ;
//            end
            begin
              rf_driver[0][11].reset()  ;
            end

//            begin
//              gen[0][12].reset()  ;
//            end
//            begin
//              drv[0][12].reset()  ;
//            end
//            begin
//              mem_check[0][12].reset()  ;
//            end
            begin
              rf_driver[0][12].reset()  ;
            end

//            begin
//              gen[0][13].reset()  ;
//            end
//            begin
//              drv[0][13].reset()  ;
//            end
//            begin
//              mem_check[0][13].reset()  ;
//            end
            begin
              rf_driver[0][13].reset()  ;
            end

//            begin
//              gen[0][14].reset()  ;
//            end
//            begin
//              drv[0][14].reset()  ;
//            end
//            begin
//              mem_check[0][14].reset()  ;
//            end
            begin
              rf_driver[0][14].reset()  ;
            end

//            begin
//              gen[0][15].reset()  ;
//            end
//            begin
//              drv[0][15].reset()  ;
//            end
//            begin
//              mem_check[0][15].reset()  ;
//            end
            begin
              rf_driver[0][15].reset()  ;
            end

//            begin
//              gen[0][16].reset()  ;
//            end
//            begin
//              drv[0][16].reset()  ;
//            end
//            begin
//              mem_check[0][16].reset()  ;
//            end
            begin
              rf_driver[0][16].reset()  ;
            end

//            begin
//              gen[0][17].reset()  ;
//            end
//            begin
//              drv[0][17].reset()  ;
//            end
//            begin
//              mem_check[0][17].reset()  ;
//            end
            begin
              rf_driver[0][17].reset()  ;
            end

//            begin
//              gen[0][18].reset()  ;
//            end
//            begin
//              drv[0][18].reset()  ;
//            end
//            begin
//              mem_check[0][18].reset()  ;
//            end
            begin
              rf_driver[0][18].reset()  ;
            end

//            begin
//              gen[0][19].reset()  ;
//            end
//            begin
//              drv[0][19].reset()  ;
//            end
//            begin
//              mem_check[0][19].reset()  ;
//            end
            begin
              rf_driver[0][19].reset()  ;
            end

//            begin
//              gen[0][20].reset()  ;
//            end
//            begin
//              drv[0][20].reset()  ;
//            end
//            begin
//              mem_check[0][20].reset()  ;
//            end
            begin
              rf_driver[0][20].reset()  ;
            end

//            begin
//              gen[0][21].reset()  ;
//            end
//            begin
//              drv[0][21].reset()  ;
//            end
//            begin
//              mem_check[0][21].reset()  ;
//            end
            begin
              rf_driver[0][21].reset()  ;
            end

//            begin
//              gen[0][22].reset()  ;
//            end
//            begin
//              drv[0][22].reset()  ;
//            end
//            begin
//              mem_check[0][22].reset()  ;
//            end
            begin
              rf_driver[0][22].reset()  ;
            end

//            begin
//              gen[0][23].reset()  ;
//            end
//            begin
//              drv[0][23].reset()  ;
//            end
//            begin
//              mem_check[0][23].reset()  ;
//            end
            begin
              rf_driver[0][23].reset()  ;
            end

//            begin
//              gen[0][24].reset()  ;
//            end
//            begin
//              drv[0][24].reset()  ;
//            end
//            begin
//              mem_check[0][24].reset()  ;
//            end
            begin
              rf_driver[0][24].reset()  ;
            end

//            begin
//              gen[0][25].reset()  ;
//            end
//            begin
//              drv[0][25].reset()  ;
//            end
//            begin
//              mem_check[0][25].reset()  ;
//            end
            begin
              rf_driver[0][25].reset()  ;
            end

//            begin
//              gen[0][26].reset()  ;
//            end
//            begin
//              drv[0][26].reset()  ;
//            end
//            begin
//              mem_check[0][26].reset()  ;
//            end
            begin
              rf_driver[0][26].reset()  ;
            end

//            begin
//              gen[0][27].reset()  ;
//            end
//            begin
//              drv[0][27].reset()  ;
//            end
//            begin
//              mem_check[0][27].reset()  ;
//            end
            begin
              rf_driver[0][27].reset()  ;
            end

//            begin
//              gen[0][28].reset()  ;
//            end
//            begin
//              drv[0][28].reset()  ;
//            end
//            begin
//              mem_check[0][28].reset()  ;
//            end
            begin
              rf_driver[0][28].reset()  ;
            end

//            begin
//              gen[0][29].reset()  ;
//            end
//            begin
//              drv[0][29].reset()  ;
//            end
//            begin
//              mem_check[0][29].reset()  ;
//            end
            begin
              rf_driver[0][29].reset()  ;
            end

//            begin
//              gen[0][30].reset()  ;
//            end
//            begin
//              drv[0][30].reset()  ;
//            end
//            begin
//              mem_check[0][30].reset()  ;
//            end
            begin
              rf_driver[0][30].reset()  ;
            end

//            begin
//              gen[0][31].reset()  ;
//            end
//            begin
//              drv[0][31].reset()  ;
//            end
//            begin
//              mem_check[0][31].reset()  ;
//            end
            begin
              rf_driver[0][31].reset()  ;
            end

//            begin
//              ldst_driver[1].reset()  ;
//            end
//            begin
//              mgr[1].reset()  ;
//            end
//            begin
//              oob_drv[1].reset()  ;
//            end
//            begin
//              up_check[1].reset()  ;
//            end
//            begin
//              gen[1][0].reset()  ;
//            end
//            begin
//              drv[1][0].reset()  ;
//            end
//            begin
//              mem_check[1][0].reset()  ;
//            end
            begin
              rf_driver[1][0].reset()  ;
            end

//            begin
//              gen[1][1].reset()  ;
//            end
//            begin
//              drv[1][1].reset()  ;
//            end
//            begin
//              mem_check[1][1].reset()  ;
//            end
            begin
              rf_driver[1][1].reset()  ;
            end

//            begin
//              gen[1][2].reset()  ;
//            end
//            begin
//              drv[1][2].reset()  ;
//            end
//            begin
//              mem_check[1][2].reset()  ;
//            end
            begin
              rf_driver[1][2].reset()  ;
            end

//            begin
//              gen[1][3].reset()  ;
//            end
//            begin
//              drv[1][3].reset()  ;
//            end
//            begin
//              mem_check[1][3].reset()  ;
//            end
            begin
              rf_driver[1][3].reset()  ;
            end

//            begin
//              gen[1][4].reset()  ;
//            end
//            begin
//              drv[1][4].reset()  ;
//            end
//            begin
//              mem_check[1][4].reset()  ;
//            end
            begin
              rf_driver[1][4].reset()  ;
            end

//            begin
//              gen[1][5].reset()  ;
//            end
//            begin
//              drv[1][5].reset()  ;
//            end
//            begin
//              mem_check[1][5].reset()  ;
//            end
            begin
              rf_driver[1][5].reset()  ;
            end

//            begin
//              gen[1][6].reset()  ;
//            end
//            begin
//              drv[1][6].reset()  ;
//            end
//            begin
//              mem_check[1][6].reset()  ;
//            end
            begin
              rf_driver[1][6].reset()  ;
            end

//            begin
//              gen[1][7].reset()  ;
//            end
//            begin
//              drv[1][7].reset()  ;
//            end
//            begin
//              mem_check[1][7].reset()  ;
//            end
            begin
              rf_driver[1][7].reset()  ;
            end

//            begin
//              gen[1][8].reset()  ;
//            end
//            begin
//              drv[1][8].reset()  ;
//            end
//            begin
//              mem_check[1][8].reset()  ;
//            end
            begin
              rf_driver[1][8].reset()  ;
            end

//            begin
//              gen[1][9].reset()  ;
//            end
//            begin
//              drv[1][9].reset()  ;
//            end
//            begin
//              mem_check[1][9].reset()  ;
//            end
            begin
              rf_driver[1][9].reset()  ;
            end

//            begin
//              gen[1][10].reset()  ;
//            end
//            begin
//              drv[1][10].reset()  ;
//            end
//            begin
//              mem_check[1][10].reset()  ;
//            end
            begin
              rf_driver[1][10].reset()  ;
            end

//            begin
//              gen[1][11].reset()  ;
//            end
//            begin
//              drv[1][11].reset()  ;
//            end
//            begin
//              mem_check[1][11].reset()  ;
//            end
            begin
              rf_driver[1][11].reset()  ;
            end

//            begin
//              gen[1][12].reset()  ;
//            end
//            begin
//              drv[1][12].reset()  ;
//            end
//            begin
//              mem_check[1][12].reset()  ;
//            end
            begin
              rf_driver[1][12].reset()  ;
            end

//            begin
//              gen[1][13].reset()  ;
//            end
//            begin
//              drv[1][13].reset()  ;
//            end
//            begin
//              mem_check[1][13].reset()  ;
//            end
            begin
              rf_driver[1][13].reset()  ;
            end

//            begin
//              gen[1][14].reset()  ;
//            end
//            begin
//              drv[1][14].reset()  ;
//            end
//            begin
//              mem_check[1][14].reset()  ;
//            end
            begin
              rf_driver[1][14].reset()  ;
            end

//            begin
//              gen[1][15].reset()  ;
//            end
//            begin
//              drv[1][15].reset()  ;
//            end
//            begin
//              mem_check[1][15].reset()  ;
//            end
            begin
              rf_driver[1][15].reset()  ;
            end

//            begin
//              gen[1][16].reset()  ;
//            end
//            begin
//              drv[1][16].reset()  ;
//            end
//            begin
//              mem_check[1][16].reset()  ;
//            end
            begin
              rf_driver[1][16].reset()  ;
            end

//            begin
//              gen[1][17].reset()  ;
//            end
//            begin
//              drv[1][17].reset()  ;
//            end
//            begin
//              mem_check[1][17].reset()  ;
//            end
            begin
              rf_driver[1][17].reset()  ;
            end

//            begin
//              gen[1][18].reset()  ;
//            end
//            begin
//              drv[1][18].reset()  ;
//            end
//            begin
//              mem_check[1][18].reset()  ;
//            end
            begin
              rf_driver[1][18].reset()  ;
            end

//            begin
//              gen[1][19].reset()  ;
//            end
//            begin
//              drv[1][19].reset()  ;
//            end
//            begin
//              mem_check[1][19].reset()  ;
//            end
            begin
              rf_driver[1][19].reset()  ;
            end

//            begin
//              gen[1][20].reset()  ;
//            end
//            begin
//              drv[1][20].reset()  ;
//            end
//            begin
//              mem_check[1][20].reset()  ;
//            end
            begin
              rf_driver[1][20].reset()  ;
            end

//            begin
//              gen[1][21].reset()  ;
//            end
//            begin
//              drv[1][21].reset()  ;
//            end
//            begin
//              mem_check[1][21].reset()  ;
//            end
            begin
              rf_driver[1][21].reset()  ;
            end

//            begin
//              gen[1][22].reset()  ;
//            end
//            begin
//              drv[1][22].reset()  ;
//            end
//            begin
//              mem_check[1][22].reset()  ;
//            end
            begin
              rf_driver[1][22].reset()  ;
            end

//            begin
//              gen[1][23].reset()  ;
//            end
//            begin
//              drv[1][23].reset()  ;
//            end
//            begin
//              mem_check[1][23].reset()  ;
//            end
            begin
              rf_driver[1][23].reset()  ;
            end

//            begin
//              gen[1][24].reset()  ;
//            end
//            begin
//              drv[1][24].reset()  ;
//            end
//            begin
//              mem_check[1][24].reset()  ;
//            end
            begin
              rf_driver[1][24].reset()  ;
            end

//            begin
//              gen[1][25].reset()  ;
//            end
//            begin
//              drv[1][25].reset()  ;
//            end
//            begin
//              mem_check[1][25].reset()  ;
//            end
            begin
              rf_driver[1][25].reset()  ;
            end

//            begin
//              gen[1][26].reset()  ;
//            end
//            begin
//              drv[1][26].reset()  ;
//            end
//            begin
//              mem_check[1][26].reset()  ;
//            end
            begin
              rf_driver[1][26].reset()  ;
            end

//            begin
//              gen[1][27].reset()  ;
//            end
//            begin
//              drv[1][27].reset()  ;
//            end
//            begin
//              mem_check[1][27].reset()  ;
//            end
            begin
              rf_driver[1][27].reset()  ;
            end

//            begin
//              gen[1][28].reset()  ;
//            end
//            begin
//              drv[1][28].reset()  ;
//            end
//            begin
//              mem_check[1][28].reset()  ;
//            end
            begin
              rf_driver[1][28].reset()  ;
            end

//            begin
//              gen[1][29].reset()  ;
//            end
//            begin
//              drv[1][29].reset()  ;
//            end
//            begin
//              mem_check[1][29].reset()  ;
//            end
            begin
              rf_driver[1][29].reset()  ;
            end

//            begin
//              gen[1][30].reset()  ;
//            end
//            begin
//              drv[1][30].reset()  ;
//            end
//            begin
//              mem_check[1][30].reset()  ;
//            end
            begin
              rf_driver[1][30].reset()  ;
            end

//            begin
//              gen[1][31].reset()  ;
//            end
//            begin
//              drv[1][31].reset()  ;
//            end
//            begin
//              mem_check[1][31].reset()  ;
//            end
            begin
              rf_driver[1][31].reset()  ;
            end

//            begin
//              ldst_driver[2].reset()  ;
//            end
//            begin
//              mgr[2].reset()  ;
//            end
//            begin
//              oob_drv[2].reset()  ;
//            end
//            begin
//              up_check[2].reset()  ;
//            end
//            begin
//              gen[2][0].reset()  ;
//            end
//            begin
//              drv[2][0].reset()  ;
//            end
//            begin
//              mem_check[2][0].reset()  ;
//            end
            begin
              rf_driver[2][0].reset()  ;
            end

//            begin
//              gen[2][1].reset()  ;
//            end
//            begin
//              drv[2][1].reset()  ;
//            end
//            begin
//              mem_check[2][1].reset()  ;
//            end
            begin
              rf_driver[2][1].reset()  ;
            end

//            begin
//              gen[2][2].reset()  ;
//            end
//            begin
//              drv[2][2].reset()  ;
//            end
//            begin
//              mem_check[2][2].reset()  ;
//            end
            begin
              rf_driver[2][2].reset()  ;
            end

//            begin
//              gen[2][3].reset()  ;
//            end
//            begin
//              drv[2][3].reset()  ;
//            end
//            begin
//              mem_check[2][3].reset()  ;
//            end
            begin
              rf_driver[2][3].reset()  ;
            end

//            begin
//              gen[2][4].reset()  ;
//            end
//            begin
//              drv[2][4].reset()  ;
//            end
//            begin
//              mem_check[2][4].reset()  ;
//            end
            begin
              rf_driver[2][4].reset()  ;
            end

//            begin
//              gen[2][5].reset()  ;
//            end
//            begin
//              drv[2][5].reset()  ;
//            end
//            begin
//              mem_check[2][5].reset()  ;
//            end
            begin
              rf_driver[2][5].reset()  ;
            end

//            begin
//              gen[2][6].reset()  ;
//            end
//            begin
//              drv[2][6].reset()  ;
//            end
//            begin
//              mem_check[2][6].reset()  ;
//            end
            begin
              rf_driver[2][6].reset()  ;
            end

//            begin
//              gen[2][7].reset()  ;
//            end
//            begin
//              drv[2][7].reset()  ;
//            end
//            begin
//              mem_check[2][7].reset()  ;
//            end
            begin
              rf_driver[2][7].reset()  ;
            end

//            begin
//              gen[2][8].reset()  ;
//            end
//            begin
//              drv[2][8].reset()  ;
//            end
//            begin
//              mem_check[2][8].reset()  ;
//            end
            begin
              rf_driver[2][8].reset()  ;
            end

//            begin
//              gen[2][9].reset()  ;
//            end
//            begin
//              drv[2][9].reset()  ;
//            end
//            begin
//              mem_check[2][9].reset()  ;
//            end
            begin
              rf_driver[2][9].reset()  ;
            end

//            begin
//              gen[2][10].reset()  ;
//            end
//            begin
//              drv[2][10].reset()  ;
//            end
//            begin
//              mem_check[2][10].reset()  ;
//            end
            begin
              rf_driver[2][10].reset()  ;
            end

//            begin
//              gen[2][11].reset()  ;
//            end
//            begin
//              drv[2][11].reset()  ;
//            end
//            begin
//              mem_check[2][11].reset()  ;
//            end
            begin
              rf_driver[2][11].reset()  ;
            end

//            begin
//              gen[2][12].reset()  ;
//            end
//            begin
//              drv[2][12].reset()  ;
//            end
//            begin
//              mem_check[2][12].reset()  ;
//            end
            begin
              rf_driver[2][12].reset()  ;
            end

//            begin
//              gen[2][13].reset()  ;
//            end
//            begin
//              drv[2][13].reset()  ;
//            end
//            begin
//              mem_check[2][13].reset()  ;
//            end
            begin
              rf_driver[2][13].reset()  ;
            end

//            begin
//              gen[2][14].reset()  ;
//            end
//            begin
//              drv[2][14].reset()  ;
//            end
//            begin
//              mem_check[2][14].reset()  ;
//            end
            begin
              rf_driver[2][14].reset()  ;
            end

//            begin
//              gen[2][15].reset()  ;
//            end
//            begin
//              drv[2][15].reset()  ;
//            end
//            begin
//              mem_check[2][15].reset()  ;
//            end
            begin
              rf_driver[2][15].reset()  ;
            end

//            begin
//              gen[2][16].reset()  ;
//            end
//            begin
//              drv[2][16].reset()  ;
//            end
//            begin
//              mem_check[2][16].reset()  ;
//            end
            begin
              rf_driver[2][16].reset()  ;
            end

//            begin
//              gen[2][17].reset()  ;
//            end
//            begin
//              drv[2][17].reset()  ;
//            end
//            begin
//              mem_check[2][17].reset()  ;
//            end
            begin
              rf_driver[2][17].reset()  ;
            end

//            begin
//              gen[2][18].reset()  ;
//            end
//            begin
//              drv[2][18].reset()  ;
//            end
//            begin
//              mem_check[2][18].reset()  ;
//            end
            begin
              rf_driver[2][18].reset()  ;
            end

//            begin
//              gen[2][19].reset()  ;
//            end
//            begin
//              drv[2][19].reset()  ;
//            end
//            begin
//              mem_check[2][19].reset()  ;
//            end
            begin
              rf_driver[2][19].reset()  ;
            end

//            begin
//              gen[2][20].reset()  ;
//            end
//            begin
//              drv[2][20].reset()  ;
//            end
//            begin
//              mem_check[2][20].reset()  ;
//            end
            begin
              rf_driver[2][20].reset()  ;
            end

//            begin
//              gen[2][21].reset()  ;
//            end
//            begin
//              drv[2][21].reset()  ;
//            end
//            begin
//              mem_check[2][21].reset()  ;
//            end
            begin
              rf_driver[2][21].reset()  ;
            end

//            begin
//              gen[2][22].reset()  ;
//            end
//            begin
//              drv[2][22].reset()  ;
//            end
//            begin
//              mem_check[2][22].reset()  ;
//            end
            begin
              rf_driver[2][22].reset()  ;
            end

//            begin
//              gen[2][23].reset()  ;
//            end
//            begin
//              drv[2][23].reset()  ;
//            end
//            begin
//              mem_check[2][23].reset()  ;
//            end
            begin
              rf_driver[2][23].reset()  ;
            end

//            begin
//              gen[2][24].reset()  ;
//            end
//            begin
//              drv[2][24].reset()  ;
//            end
//            begin
//              mem_check[2][24].reset()  ;
//            end
            begin
              rf_driver[2][24].reset()  ;
            end

//            begin
//              gen[2][25].reset()  ;
//            end
//            begin
//              drv[2][25].reset()  ;
//            end
//            begin
//              mem_check[2][25].reset()  ;
//            end
            begin
              rf_driver[2][25].reset()  ;
            end

//            begin
//              gen[2][26].reset()  ;
//            end
//            begin
//              drv[2][26].reset()  ;
//            end
//            begin
//              mem_check[2][26].reset()  ;
//            end
            begin
              rf_driver[2][26].reset()  ;
            end

//            begin
//              gen[2][27].reset()  ;
//            end
//            begin
//              drv[2][27].reset()  ;
//            end
//            begin
//              mem_check[2][27].reset()  ;
//            end
            begin
              rf_driver[2][27].reset()  ;
            end

//            begin
//              gen[2][28].reset()  ;
//            end
//            begin
//              drv[2][28].reset()  ;
//            end
//            begin
//              mem_check[2][28].reset()  ;
//            end
            begin
              rf_driver[2][28].reset()  ;
            end

//            begin
//              gen[2][29].reset()  ;
//            end
//            begin
//              drv[2][29].reset()  ;
//            end
//            begin
//              mem_check[2][29].reset()  ;
//            end
            begin
              rf_driver[2][29].reset()  ;
            end

//            begin
//              gen[2][30].reset()  ;
//            end
//            begin
//              drv[2][30].reset()  ;
//            end
//            begin
//              mem_check[2][30].reset()  ;
//            end
            begin
              rf_driver[2][30].reset()  ;
            end

//            begin
//              gen[2][31].reset()  ;
//            end
//            begin
//              drv[2][31].reset()  ;
//            end
//            begin
//              mem_check[2][31].reset()  ;
//            end
            begin
              rf_driver[2][31].reset()  ;
            end

//            begin
//              ldst_driver[3].reset()  ;
//            end
//            begin
//              mgr[3].reset()  ;
//            end
//            begin
//              oob_drv[3].reset()  ;
//            end
//            begin
//              up_check[3].reset()  ;
//            end
//            begin
//              gen[3][0].reset()  ;
//            end
//            begin
//              drv[3][0].reset()  ;
//            end
//            begin
//              mem_check[3][0].reset()  ;
//            end
            begin
              rf_driver[3][0].reset()  ;
            end

//            begin
//              gen[3][1].reset()  ;
//            end
//            begin
//              drv[3][1].reset()  ;
//            end
//            begin
//              mem_check[3][1].reset()  ;
//            end
            begin
              rf_driver[3][1].reset()  ;
            end

//            begin
//              gen[3][2].reset()  ;
//            end
//            begin
//              drv[3][2].reset()  ;
//            end
//            begin
//              mem_check[3][2].reset()  ;
//            end
            begin
              rf_driver[3][2].reset()  ;
            end

//            begin
//              gen[3][3].reset()  ;
//            end
//            begin
//              drv[3][3].reset()  ;
//            end
//            begin
//              mem_check[3][3].reset()  ;
//            end
            begin
              rf_driver[3][3].reset()  ;
            end

//            begin
//              gen[3][4].reset()  ;
//            end
//            begin
//              drv[3][4].reset()  ;
//            end
//            begin
//              mem_check[3][4].reset()  ;
//            end
            begin
              rf_driver[3][4].reset()  ;
            end

//            begin
//              gen[3][5].reset()  ;
//            end
//            begin
//              drv[3][5].reset()  ;
//            end
//            begin
//              mem_check[3][5].reset()  ;
//            end
            begin
              rf_driver[3][5].reset()  ;
            end

//            begin
//              gen[3][6].reset()  ;
//            end
//            begin
//              drv[3][6].reset()  ;
//            end
//            begin
//              mem_check[3][6].reset()  ;
//            end
            begin
              rf_driver[3][6].reset()  ;
            end

//            begin
//              gen[3][7].reset()  ;
//            end
//            begin
//              drv[3][7].reset()  ;
//            end
//            begin
//              mem_check[3][7].reset()  ;
//            end
            begin
              rf_driver[3][7].reset()  ;
            end

//            begin
//              gen[3][8].reset()  ;
//            end
//            begin
//              drv[3][8].reset()  ;
//            end
//            begin
//              mem_check[3][8].reset()  ;
//            end
            begin
              rf_driver[3][8].reset()  ;
            end

//            begin
//              gen[3][9].reset()  ;
//            end
//            begin
//              drv[3][9].reset()  ;
//            end
//            begin
//              mem_check[3][9].reset()  ;
//            end
            begin
              rf_driver[3][9].reset()  ;
            end

//            begin
//              gen[3][10].reset()  ;
//            end
//            begin
//              drv[3][10].reset()  ;
//            end
//            begin
//              mem_check[3][10].reset()  ;
//            end
            begin
              rf_driver[3][10].reset()  ;
            end

//            begin
//              gen[3][11].reset()  ;
//            end
//            begin
//              drv[3][11].reset()  ;
//            end
//            begin
//              mem_check[3][11].reset()  ;
//            end
            begin
              rf_driver[3][11].reset()  ;
            end

//            begin
//              gen[3][12].reset()  ;
//            end
//            begin
//              drv[3][12].reset()  ;
//            end
//            begin
//              mem_check[3][12].reset()  ;
//            end
            begin
              rf_driver[3][12].reset()  ;
            end

//            begin
//              gen[3][13].reset()  ;
//            end
//            begin
//              drv[3][13].reset()  ;
//            end
//            begin
//              mem_check[3][13].reset()  ;
//            end
            begin
              rf_driver[3][13].reset()  ;
            end

//            begin
//              gen[3][14].reset()  ;
//            end
//            begin
//              drv[3][14].reset()  ;
//            end
//            begin
//              mem_check[3][14].reset()  ;
//            end
            begin
              rf_driver[3][14].reset()  ;
            end

//            begin
//              gen[3][15].reset()  ;
//            end
//            begin
//              drv[3][15].reset()  ;
//            end
//            begin
//              mem_check[3][15].reset()  ;
//            end
            begin
              rf_driver[3][15].reset()  ;
            end

//            begin
//              gen[3][16].reset()  ;
//            end
//            begin
//              drv[3][16].reset()  ;
//            end
//            begin
//              mem_check[3][16].reset()  ;
//            end
            begin
              rf_driver[3][16].reset()  ;
            end

//            begin
//              gen[3][17].reset()  ;
//            end
//            begin
//              drv[3][17].reset()  ;
//            end
//            begin
//              mem_check[3][17].reset()  ;
//            end
            begin
              rf_driver[3][17].reset()  ;
            end

//            begin
//              gen[3][18].reset()  ;
//            end
//            begin
//              drv[3][18].reset()  ;
//            end
//            begin
//              mem_check[3][18].reset()  ;
//            end
            begin
              rf_driver[3][18].reset()  ;
            end

//            begin
//              gen[3][19].reset()  ;
//            end
//            begin
//              drv[3][19].reset()  ;
//            end
//            begin
//              mem_check[3][19].reset()  ;
//            end
            begin
              rf_driver[3][19].reset()  ;
            end

//            begin
//              gen[3][20].reset()  ;
//            end
//            begin
//              drv[3][20].reset()  ;
//            end
//            begin
//              mem_check[3][20].reset()  ;
//            end
            begin
              rf_driver[3][20].reset()  ;
            end

//            begin
//              gen[3][21].reset()  ;
//            end
//            begin
//              drv[3][21].reset()  ;
//            end
//            begin
//              mem_check[3][21].reset()  ;
//            end
            begin
              rf_driver[3][21].reset()  ;
            end

//            begin
//              gen[3][22].reset()  ;
//            end
//            begin
//              drv[3][22].reset()  ;
//            end
//            begin
//              mem_check[3][22].reset()  ;
//            end
            begin
              rf_driver[3][22].reset()  ;
            end

//            begin
//              gen[3][23].reset()  ;
//            end
//            begin
//              drv[3][23].reset()  ;
//            end
//            begin
//              mem_check[3][23].reset()  ;
//            end
            begin
              rf_driver[3][23].reset()  ;
            end

//            begin
//              gen[3][24].reset()  ;
//            end
//            begin
//              drv[3][24].reset()  ;
//            end
//            begin
//              mem_check[3][24].reset()  ;
//            end
            begin
              rf_driver[3][24].reset()  ;
            end

//            begin
//              gen[3][25].reset()  ;
//            end
//            begin
//              drv[3][25].reset()  ;
//            end
//            begin
//              mem_check[3][25].reset()  ;
//            end
            begin
              rf_driver[3][25].reset()  ;
            end

//            begin
//              gen[3][26].reset()  ;
//            end
//            begin
//              drv[3][26].reset()  ;
//            end
//            begin
//              mem_check[3][26].reset()  ;
//            end
            begin
              rf_driver[3][26].reset()  ;
            end

//            begin
//              gen[3][27].reset()  ;
//            end
//            begin
//              drv[3][27].reset()  ;
//            end
//            begin
//              mem_check[3][27].reset()  ;
//            end
            begin
              rf_driver[3][27].reset()  ;
            end

//            begin
//              gen[3][28].reset()  ;
//            end
//            begin
//              drv[3][28].reset()  ;
//            end
//            begin
//              mem_check[3][28].reset()  ;
//            end
            begin
              rf_driver[3][28].reset()  ;
            end

//            begin
//              gen[3][29].reset()  ;
//            end
//            begin
//              drv[3][29].reset()  ;
//            end
//            begin
//              mem_check[3][29].reset()  ;
//            end
            begin
              rf_driver[3][29].reset()  ;
            end

//            begin
//              gen[3][30].reset()  ;
//            end
//            begin
//              drv[3][30].reset()  ;
//            end
//            begin
//              mem_check[3][30].reset()  ;
//            end
            begin
              rf_driver[3][30].reset()  ;
            end

//            begin
//              gen[3][31].reset()  ;
//            end
//            begin
//              drv[3][31].reset()  ;
//            end
//            begin
//              mem_check[3][31].reset()  ;
//            end
            begin
              rf_driver[3][31].reset()  ;
            end
