
  assign   pe0__stu__valid                =  pe_inst[0].pe__stu__valid     ;
  assign   pe0__stu__cntl                 =  pe_inst[0].pe__stu__cntl      ;
  assign   pe_inst[0].stu__pe__ready      =  stu__pe0__ready               ;
  assign   pe0__stu__type                 =  pe_inst[0].pe__stu__type      ;
  assign   pe0__stu__data                 =  pe_inst[0].pe__stu__data      ;
  assign   pe0__stu__oob_data             =  pe_inst[0].pe__stu__oob_data  ;

  assign   pe1__stu__valid                =  pe_inst[1].pe__stu__valid     ;
  assign   pe1__stu__cntl                 =  pe_inst[1].pe__stu__cntl      ;
  assign   pe_inst[1].stu__pe__ready      =  stu__pe1__ready               ;
  assign   pe1__stu__type                 =  pe_inst[1].pe__stu__type      ;
  assign   pe1__stu__data                 =  pe_inst[1].pe__stu__data      ;
  assign   pe1__stu__oob_data             =  pe_inst[1].pe__stu__oob_data  ;

  assign   pe2__stu__valid                =  pe_inst[2].pe__stu__valid     ;
  assign   pe2__stu__cntl                 =  pe_inst[2].pe__stu__cntl      ;
  assign   pe_inst[2].stu__pe__ready      =  stu__pe2__ready               ;
  assign   pe2__stu__type                 =  pe_inst[2].pe__stu__type      ;
  assign   pe2__stu__data                 =  pe_inst[2].pe__stu__data      ;
  assign   pe2__stu__oob_data             =  pe_inst[2].pe__stu__oob_data  ;

  assign   pe3__stu__valid                =  pe_inst[3].pe__stu__valid     ;
  assign   pe3__stu__cntl                 =  pe_inst[3].pe__stu__cntl      ;
  assign   pe_inst[3].stu__pe__ready      =  stu__pe3__ready               ;
  assign   pe3__stu__type                 =  pe_inst[3].pe__stu__type      ;
  assign   pe3__stu__data                 =  pe_inst[3].pe__stu__data      ;
  assign   pe3__stu__oob_data             =  pe_inst[3].pe__stu__oob_data  ;

  assign   pe4__stu__valid                =  pe_inst[4].pe__stu__valid     ;
  assign   pe4__stu__cntl                 =  pe_inst[4].pe__stu__cntl      ;
  assign   pe_inst[4].stu__pe__ready      =  stu__pe4__ready               ;
  assign   pe4__stu__type                 =  pe_inst[4].pe__stu__type      ;
  assign   pe4__stu__data                 =  pe_inst[4].pe__stu__data      ;
  assign   pe4__stu__oob_data             =  pe_inst[4].pe__stu__oob_data  ;

  assign   pe5__stu__valid                =  pe_inst[5].pe__stu__valid     ;
  assign   pe5__stu__cntl                 =  pe_inst[5].pe__stu__cntl      ;
  assign   pe_inst[5].stu__pe__ready      =  stu__pe5__ready               ;
  assign   pe5__stu__type                 =  pe_inst[5].pe__stu__type      ;
  assign   pe5__stu__data                 =  pe_inst[5].pe__stu__data      ;
  assign   pe5__stu__oob_data             =  pe_inst[5].pe__stu__oob_data  ;

  assign   pe6__stu__valid                =  pe_inst[6].pe__stu__valid     ;
  assign   pe6__stu__cntl                 =  pe_inst[6].pe__stu__cntl      ;
  assign   pe_inst[6].stu__pe__ready      =  stu__pe6__ready               ;
  assign   pe6__stu__type                 =  pe_inst[6].pe__stu__type      ;
  assign   pe6__stu__data                 =  pe_inst[6].pe__stu__data      ;
  assign   pe6__stu__oob_data             =  pe_inst[6].pe__stu__oob_data  ;

  assign   pe7__stu__valid                =  pe_inst[7].pe__stu__valid     ;
  assign   pe7__stu__cntl                 =  pe_inst[7].pe__stu__cntl      ;
  assign   pe_inst[7].stu__pe__ready      =  stu__pe7__ready               ;
  assign   pe7__stu__type                 =  pe_inst[7].pe__stu__type      ;
  assign   pe7__stu__data                 =  pe_inst[7].pe__stu__data      ;
  assign   pe7__stu__oob_data             =  pe_inst[7].pe__stu__oob_data  ;

  assign   pe8__stu__valid                =  pe_inst[8].pe__stu__valid     ;
  assign   pe8__stu__cntl                 =  pe_inst[8].pe__stu__cntl      ;
  assign   pe_inst[8].stu__pe__ready      =  stu__pe8__ready               ;
  assign   pe8__stu__type                 =  pe_inst[8].pe__stu__type      ;
  assign   pe8__stu__data                 =  pe_inst[8].pe__stu__data      ;
  assign   pe8__stu__oob_data             =  pe_inst[8].pe__stu__oob_data  ;

  assign   pe9__stu__valid                =  pe_inst[9].pe__stu__valid     ;
  assign   pe9__stu__cntl                 =  pe_inst[9].pe__stu__cntl      ;
  assign   pe_inst[9].stu__pe__ready      =  stu__pe9__ready               ;
  assign   pe9__stu__type                 =  pe_inst[9].pe__stu__type      ;
  assign   pe9__stu__data                 =  pe_inst[9].pe__stu__data      ;
  assign   pe9__stu__oob_data             =  pe_inst[9].pe__stu__oob_data  ;

  assign   pe10__stu__valid                =  pe_inst[10].pe__stu__valid     ;
  assign   pe10__stu__cntl                 =  pe_inst[10].pe__stu__cntl      ;
  assign   pe_inst[10].stu__pe__ready      =  stu__pe10__ready               ;
  assign   pe10__stu__type                 =  pe_inst[10].pe__stu__type      ;
  assign   pe10__stu__data                 =  pe_inst[10].pe__stu__data      ;
  assign   pe10__stu__oob_data             =  pe_inst[10].pe__stu__oob_data  ;

  assign   pe11__stu__valid                =  pe_inst[11].pe__stu__valid     ;
  assign   pe11__stu__cntl                 =  pe_inst[11].pe__stu__cntl      ;
  assign   pe_inst[11].stu__pe__ready      =  stu__pe11__ready               ;
  assign   pe11__stu__type                 =  pe_inst[11].pe__stu__type      ;
  assign   pe11__stu__data                 =  pe_inst[11].pe__stu__data      ;
  assign   pe11__stu__oob_data             =  pe_inst[11].pe__stu__oob_data  ;

  assign   pe12__stu__valid                =  pe_inst[12].pe__stu__valid     ;
  assign   pe12__stu__cntl                 =  pe_inst[12].pe__stu__cntl      ;
  assign   pe_inst[12].stu__pe__ready      =  stu__pe12__ready               ;
  assign   pe12__stu__type                 =  pe_inst[12].pe__stu__type      ;
  assign   pe12__stu__data                 =  pe_inst[12].pe__stu__data      ;
  assign   pe12__stu__oob_data             =  pe_inst[12].pe__stu__oob_data  ;

  assign   pe13__stu__valid                =  pe_inst[13].pe__stu__valid     ;
  assign   pe13__stu__cntl                 =  pe_inst[13].pe__stu__cntl      ;
  assign   pe_inst[13].stu__pe__ready      =  stu__pe13__ready               ;
  assign   pe13__stu__type                 =  pe_inst[13].pe__stu__type      ;
  assign   pe13__stu__data                 =  pe_inst[13].pe__stu__data      ;
  assign   pe13__stu__oob_data             =  pe_inst[13].pe__stu__oob_data  ;

  assign   pe14__stu__valid                =  pe_inst[14].pe__stu__valid     ;
  assign   pe14__stu__cntl                 =  pe_inst[14].pe__stu__cntl      ;
  assign   pe_inst[14].stu__pe__ready      =  stu__pe14__ready               ;
  assign   pe14__stu__type                 =  pe_inst[14].pe__stu__type      ;
  assign   pe14__stu__data                 =  pe_inst[14].pe__stu__data      ;
  assign   pe14__stu__oob_data             =  pe_inst[14].pe__stu__oob_data  ;

  assign   pe15__stu__valid                =  pe_inst[15].pe__stu__valid     ;
  assign   pe15__stu__cntl                 =  pe_inst[15].pe__stu__cntl      ;
  assign   pe_inst[15].stu__pe__ready      =  stu__pe15__ready               ;
  assign   pe15__stu__type                 =  pe_inst[15].pe__stu__type      ;
  assign   pe15__stu__data                 =  pe_inst[15].pe__stu__data      ;
  assign   pe15__stu__oob_data             =  pe_inst[15].pe__stu__oob_data  ;

  assign   pe16__stu__valid                =  pe_inst[16].pe__stu__valid     ;
  assign   pe16__stu__cntl                 =  pe_inst[16].pe__stu__cntl      ;
  assign   pe_inst[16].stu__pe__ready      =  stu__pe16__ready               ;
  assign   pe16__stu__type                 =  pe_inst[16].pe__stu__type      ;
  assign   pe16__stu__data                 =  pe_inst[16].pe__stu__data      ;
  assign   pe16__stu__oob_data             =  pe_inst[16].pe__stu__oob_data  ;

  assign   pe17__stu__valid                =  pe_inst[17].pe__stu__valid     ;
  assign   pe17__stu__cntl                 =  pe_inst[17].pe__stu__cntl      ;
  assign   pe_inst[17].stu__pe__ready      =  stu__pe17__ready               ;
  assign   pe17__stu__type                 =  pe_inst[17].pe__stu__type      ;
  assign   pe17__stu__data                 =  pe_inst[17].pe__stu__data      ;
  assign   pe17__stu__oob_data             =  pe_inst[17].pe__stu__oob_data  ;

  assign   pe18__stu__valid                =  pe_inst[18].pe__stu__valid     ;
  assign   pe18__stu__cntl                 =  pe_inst[18].pe__stu__cntl      ;
  assign   pe_inst[18].stu__pe__ready      =  stu__pe18__ready               ;
  assign   pe18__stu__type                 =  pe_inst[18].pe__stu__type      ;
  assign   pe18__stu__data                 =  pe_inst[18].pe__stu__data      ;
  assign   pe18__stu__oob_data             =  pe_inst[18].pe__stu__oob_data  ;

  assign   pe19__stu__valid                =  pe_inst[19].pe__stu__valid     ;
  assign   pe19__stu__cntl                 =  pe_inst[19].pe__stu__cntl      ;
  assign   pe_inst[19].stu__pe__ready      =  stu__pe19__ready               ;
  assign   pe19__stu__type                 =  pe_inst[19].pe__stu__type      ;
  assign   pe19__stu__data                 =  pe_inst[19].pe__stu__data      ;
  assign   pe19__stu__oob_data             =  pe_inst[19].pe__stu__oob_data  ;

  assign   pe20__stu__valid                =  pe_inst[20].pe__stu__valid     ;
  assign   pe20__stu__cntl                 =  pe_inst[20].pe__stu__cntl      ;
  assign   pe_inst[20].stu__pe__ready      =  stu__pe20__ready               ;
  assign   pe20__stu__type                 =  pe_inst[20].pe__stu__type      ;
  assign   pe20__stu__data                 =  pe_inst[20].pe__stu__data      ;
  assign   pe20__stu__oob_data             =  pe_inst[20].pe__stu__oob_data  ;

  assign   pe21__stu__valid                =  pe_inst[21].pe__stu__valid     ;
  assign   pe21__stu__cntl                 =  pe_inst[21].pe__stu__cntl      ;
  assign   pe_inst[21].stu__pe__ready      =  stu__pe21__ready               ;
  assign   pe21__stu__type                 =  pe_inst[21].pe__stu__type      ;
  assign   pe21__stu__data                 =  pe_inst[21].pe__stu__data      ;
  assign   pe21__stu__oob_data             =  pe_inst[21].pe__stu__oob_data  ;

  assign   pe22__stu__valid                =  pe_inst[22].pe__stu__valid     ;
  assign   pe22__stu__cntl                 =  pe_inst[22].pe__stu__cntl      ;
  assign   pe_inst[22].stu__pe__ready      =  stu__pe22__ready               ;
  assign   pe22__stu__type                 =  pe_inst[22].pe__stu__type      ;
  assign   pe22__stu__data                 =  pe_inst[22].pe__stu__data      ;
  assign   pe22__stu__oob_data             =  pe_inst[22].pe__stu__oob_data  ;

  assign   pe23__stu__valid                =  pe_inst[23].pe__stu__valid     ;
  assign   pe23__stu__cntl                 =  pe_inst[23].pe__stu__cntl      ;
  assign   pe_inst[23].stu__pe__ready      =  stu__pe23__ready               ;
  assign   pe23__stu__type                 =  pe_inst[23].pe__stu__type      ;
  assign   pe23__stu__data                 =  pe_inst[23].pe__stu__data      ;
  assign   pe23__stu__oob_data             =  pe_inst[23].pe__stu__oob_data  ;

  assign   pe24__stu__valid                =  pe_inst[24].pe__stu__valid     ;
  assign   pe24__stu__cntl                 =  pe_inst[24].pe__stu__cntl      ;
  assign   pe_inst[24].stu__pe__ready      =  stu__pe24__ready               ;
  assign   pe24__stu__type                 =  pe_inst[24].pe__stu__type      ;
  assign   pe24__stu__data                 =  pe_inst[24].pe__stu__data      ;
  assign   pe24__stu__oob_data             =  pe_inst[24].pe__stu__oob_data  ;

  assign   pe25__stu__valid                =  pe_inst[25].pe__stu__valid     ;
  assign   pe25__stu__cntl                 =  pe_inst[25].pe__stu__cntl      ;
  assign   pe_inst[25].stu__pe__ready      =  stu__pe25__ready               ;
  assign   pe25__stu__type                 =  pe_inst[25].pe__stu__type      ;
  assign   pe25__stu__data                 =  pe_inst[25].pe__stu__data      ;
  assign   pe25__stu__oob_data             =  pe_inst[25].pe__stu__oob_data  ;

  assign   pe26__stu__valid                =  pe_inst[26].pe__stu__valid     ;
  assign   pe26__stu__cntl                 =  pe_inst[26].pe__stu__cntl      ;
  assign   pe_inst[26].stu__pe__ready      =  stu__pe26__ready               ;
  assign   pe26__stu__type                 =  pe_inst[26].pe__stu__type      ;
  assign   pe26__stu__data                 =  pe_inst[26].pe__stu__data      ;
  assign   pe26__stu__oob_data             =  pe_inst[26].pe__stu__oob_data  ;

  assign   pe27__stu__valid                =  pe_inst[27].pe__stu__valid     ;
  assign   pe27__stu__cntl                 =  pe_inst[27].pe__stu__cntl      ;
  assign   pe_inst[27].stu__pe__ready      =  stu__pe27__ready               ;
  assign   pe27__stu__type                 =  pe_inst[27].pe__stu__type      ;
  assign   pe27__stu__data                 =  pe_inst[27].pe__stu__data      ;
  assign   pe27__stu__oob_data             =  pe_inst[27].pe__stu__oob_data  ;

  assign   pe28__stu__valid                =  pe_inst[28].pe__stu__valid     ;
  assign   pe28__stu__cntl                 =  pe_inst[28].pe__stu__cntl      ;
  assign   pe_inst[28].stu__pe__ready      =  stu__pe28__ready               ;
  assign   pe28__stu__type                 =  pe_inst[28].pe__stu__type      ;
  assign   pe28__stu__data                 =  pe_inst[28].pe__stu__data      ;
  assign   pe28__stu__oob_data             =  pe_inst[28].pe__stu__oob_data  ;

  assign   pe29__stu__valid                =  pe_inst[29].pe__stu__valid     ;
  assign   pe29__stu__cntl                 =  pe_inst[29].pe__stu__cntl      ;
  assign   pe_inst[29].stu__pe__ready      =  stu__pe29__ready               ;
  assign   pe29__stu__type                 =  pe_inst[29].pe__stu__type      ;
  assign   pe29__stu__data                 =  pe_inst[29].pe__stu__data      ;
  assign   pe29__stu__oob_data             =  pe_inst[29].pe__stu__oob_data  ;

  assign   pe30__stu__valid                =  pe_inst[30].pe__stu__valid     ;
  assign   pe30__stu__cntl                 =  pe_inst[30].pe__stu__cntl      ;
  assign   pe_inst[30].stu__pe__ready      =  stu__pe30__ready               ;
  assign   pe30__stu__type                 =  pe_inst[30].pe__stu__type      ;
  assign   pe30__stu__data                 =  pe_inst[30].pe__stu__data      ;
  assign   pe30__stu__oob_data             =  pe_inst[30].pe__stu__oob_data  ;

  assign   pe31__stu__valid                =  pe_inst[31].pe__stu__valid     ;
  assign   pe31__stu__cntl                 =  pe_inst[31].pe__stu__cntl      ;
  assign   pe_inst[31].stu__pe__ready      =  stu__pe31__ready               ;
  assign   pe31__stu__type                 =  pe_inst[31].pe__stu__type      ;
  assign   pe31__stu__data                 =  pe_inst[31].pe__stu__data      ;
  assign   pe31__stu__oob_data             =  pe_inst[31].pe__stu__oob_data  ;

  assign   pe32__stu__valid                =  pe_inst[32].pe__stu__valid     ;
  assign   pe32__stu__cntl                 =  pe_inst[32].pe__stu__cntl      ;
  assign   pe_inst[32].stu__pe__ready      =  stu__pe32__ready               ;
  assign   pe32__stu__type                 =  pe_inst[32].pe__stu__type      ;
  assign   pe32__stu__data                 =  pe_inst[32].pe__stu__data      ;
  assign   pe32__stu__oob_data             =  pe_inst[32].pe__stu__oob_data  ;

  assign   pe33__stu__valid                =  pe_inst[33].pe__stu__valid     ;
  assign   pe33__stu__cntl                 =  pe_inst[33].pe__stu__cntl      ;
  assign   pe_inst[33].stu__pe__ready      =  stu__pe33__ready               ;
  assign   pe33__stu__type                 =  pe_inst[33].pe__stu__type      ;
  assign   pe33__stu__data                 =  pe_inst[33].pe__stu__data      ;
  assign   pe33__stu__oob_data             =  pe_inst[33].pe__stu__oob_data  ;

  assign   pe34__stu__valid                =  pe_inst[34].pe__stu__valid     ;
  assign   pe34__stu__cntl                 =  pe_inst[34].pe__stu__cntl      ;
  assign   pe_inst[34].stu__pe__ready      =  stu__pe34__ready               ;
  assign   pe34__stu__type                 =  pe_inst[34].pe__stu__type      ;
  assign   pe34__stu__data                 =  pe_inst[34].pe__stu__data      ;
  assign   pe34__stu__oob_data             =  pe_inst[34].pe__stu__oob_data  ;

  assign   pe35__stu__valid                =  pe_inst[35].pe__stu__valid     ;
  assign   pe35__stu__cntl                 =  pe_inst[35].pe__stu__cntl      ;
  assign   pe_inst[35].stu__pe__ready      =  stu__pe35__ready               ;
  assign   pe35__stu__type                 =  pe_inst[35].pe__stu__type      ;
  assign   pe35__stu__data                 =  pe_inst[35].pe__stu__data      ;
  assign   pe35__stu__oob_data             =  pe_inst[35].pe__stu__oob_data  ;

  assign   pe36__stu__valid                =  pe_inst[36].pe__stu__valid     ;
  assign   pe36__stu__cntl                 =  pe_inst[36].pe__stu__cntl      ;
  assign   pe_inst[36].stu__pe__ready      =  stu__pe36__ready               ;
  assign   pe36__stu__type                 =  pe_inst[36].pe__stu__type      ;
  assign   pe36__stu__data                 =  pe_inst[36].pe__stu__data      ;
  assign   pe36__stu__oob_data             =  pe_inst[36].pe__stu__oob_data  ;

  assign   pe37__stu__valid                =  pe_inst[37].pe__stu__valid     ;
  assign   pe37__stu__cntl                 =  pe_inst[37].pe__stu__cntl      ;
  assign   pe_inst[37].stu__pe__ready      =  stu__pe37__ready               ;
  assign   pe37__stu__type                 =  pe_inst[37].pe__stu__type      ;
  assign   pe37__stu__data                 =  pe_inst[37].pe__stu__data      ;
  assign   pe37__stu__oob_data             =  pe_inst[37].pe__stu__oob_data  ;

  assign   pe38__stu__valid                =  pe_inst[38].pe__stu__valid     ;
  assign   pe38__stu__cntl                 =  pe_inst[38].pe__stu__cntl      ;
  assign   pe_inst[38].stu__pe__ready      =  stu__pe38__ready               ;
  assign   pe38__stu__type                 =  pe_inst[38].pe__stu__type      ;
  assign   pe38__stu__data                 =  pe_inst[38].pe__stu__data      ;
  assign   pe38__stu__oob_data             =  pe_inst[38].pe__stu__oob_data  ;

  assign   pe39__stu__valid                =  pe_inst[39].pe__stu__valid     ;
  assign   pe39__stu__cntl                 =  pe_inst[39].pe__stu__cntl      ;
  assign   pe_inst[39].stu__pe__ready      =  stu__pe39__ready               ;
  assign   pe39__stu__type                 =  pe_inst[39].pe__stu__type      ;
  assign   pe39__stu__data                 =  pe_inst[39].pe__stu__data      ;
  assign   pe39__stu__oob_data             =  pe_inst[39].pe__stu__oob_data  ;

  assign   pe40__stu__valid                =  pe_inst[40].pe__stu__valid     ;
  assign   pe40__stu__cntl                 =  pe_inst[40].pe__stu__cntl      ;
  assign   pe_inst[40].stu__pe__ready      =  stu__pe40__ready               ;
  assign   pe40__stu__type                 =  pe_inst[40].pe__stu__type      ;
  assign   pe40__stu__data                 =  pe_inst[40].pe__stu__data      ;
  assign   pe40__stu__oob_data             =  pe_inst[40].pe__stu__oob_data  ;

  assign   pe41__stu__valid                =  pe_inst[41].pe__stu__valid     ;
  assign   pe41__stu__cntl                 =  pe_inst[41].pe__stu__cntl      ;
  assign   pe_inst[41].stu__pe__ready      =  stu__pe41__ready               ;
  assign   pe41__stu__type                 =  pe_inst[41].pe__stu__type      ;
  assign   pe41__stu__data                 =  pe_inst[41].pe__stu__data      ;
  assign   pe41__stu__oob_data             =  pe_inst[41].pe__stu__oob_data  ;

  assign   pe42__stu__valid                =  pe_inst[42].pe__stu__valid     ;
  assign   pe42__stu__cntl                 =  pe_inst[42].pe__stu__cntl      ;
  assign   pe_inst[42].stu__pe__ready      =  stu__pe42__ready               ;
  assign   pe42__stu__type                 =  pe_inst[42].pe__stu__type      ;
  assign   pe42__stu__data                 =  pe_inst[42].pe__stu__data      ;
  assign   pe42__stu__oob_data             =  pe_inst[42].pe__stu__oob_data  ;

  assign   pe43__stu__valid                =  pe_inst[43].pe__stu__valid     ;
  assign   pe43__stu__cntl                 =  pe_inst[43].pe__stu__cntl      ;
  assign   pe_inst[43].stu__pe__ready      =  stu__pe43__ready               ;
  assign   pe43__stu__type                 =  pe_inst[43].pe__stu__type      ;
  assign   pe43__stu__data                 =  pe_inst[43].pe__stu__data      ;
  assign   pe43__stu__oob_data             =  pe_inst[43].pe__stu__oob_data  ;

  assign   pe44__stu__valid                =  pe_inst[44].pe__stu__valid     ;
  assign   pe44__stu__cntl                 =  pe_inst[44].pe__stu__cntl      ;
  assign   pe_inst[44].stu__pe__ready      =  stu__pe44__ready               ;
  assign   pe44__stu__type                 =  pe_inst[44].pe__stu__type      ;
  assign   pe44__stu__data                 =  pe_inst[44].pe__stu__data      ;
  assign   pe44__stu__oob_data             =  pe_inst[44].pe__stu__oob_data  ;

  assign   pe45__stu__valid                =  pe_inst[45].pe__stu__valid     ;
  assign   pe45__stu__cntl                 =  pe_inst[45].pe__stu__cntl      ;
  assign   pe_inst[45].stu__pe__ready      =  stu__pe45__ready               ;
  assign   pe45__stu__type                 =  pe_inst[45].pe__stu__type      ;
  assign   pe45__stu__data                 =  pe_inst[45].pe__stu__data      ;
  assign   pe45__stu__oob_data             =  pe_inst[45].pe__stu__oob_data  ;

  assign   pe46__stu__valid                =  pe_inst[46].pe__stu__valid     ;
  assign   pe46__stu__cntl                 =  pe_inst[46].pe__stu__cntl      ;
  assign   pe_inst[46].stu__pe__ready      =  stu__pe46__ready               ;
  assign   pe46__stu__type                 =  pe_inst[46].pe__stu__type      ;
  assign   pe46__stu__data                 =  pe_inst[46].pe__stu__data      ;
  assign   pe46__stu__oob_data             =  pe_inst[46].pe__stu__oob_data  ;

  assign   pe47__stu__valid                =  pe_inst[47].pe__stu__valid     ;
  assign   pe47__stu__cntl                 =  pe_inst[47].pe__stu__cntl      ;
  assign   pe_inst[47].stu__pe__ready      =  stu__pe47__ready               ;
  assign   pe47__stu__type                 =  pe_inst[47].pe__stu__type      ;
  assign   pe47__stu__data                 =  pe_inst[47].pe__stu__data      ;
  assign   pe47__stu__oob_data             =  pe_inst[47].pe__stu__oob_data  ;

  assign   pe48__stu__valid                =  pe_inst[48].pe__stu__valid     ;
  assign   pe48__stu__cntl                 =  pe_inst[48].pe__stu__cntl      ;
  assign   pe_inst[48].stu__pe__ready      =  stu__pe48__ready               ;
  assign   pe48__stu__type                 =  pe_inst[48].pe__stu__type      ;
  assign   pe48__stu__data                 =  pe_inst[48].pe__stu__data      ;
  assign   pe48__stu__oob_data             =  pe_inst[48].pe__stu__oob_data  ;

  assign   pe49__stu__valid                =  pe_inst[49].pe__stu__valid     ;
  assign   pe49__stu__cntl                 =  pe_inst[49].pe__stu__cntl      ;
  assign   pe_inst[49].stu__pe__ready      =  stu__pe49__ready               ;
  assign   pe49__stu__type                 =  pe_inst[49].pe__stu__type      ;
  assign   pe49__stu__data                 =  pe_inst[49].pe__stu__data      ;
  assign   pe49__stu__oob_data             =  pe_inst[49].pe__stu__oob_data  ;

  assign   pe50__stu__valid                =  pe_inst[50].pe__stu__valid     ;
  assign   pe50__stu__cntl                 =  pe_inst[50].pe__stu__cntl      ;
  assign   pe_inst[50].stu__pe__ready      =  stu__pe50__ready               ;
  assign   pe50__stu__type                 =  pe_inst[50].pe__stu__type      ;
  assign   pe50__stu__data                 =  pe_inst[50].pe__stu__data      ;
  assign   pe50__stu__oob_data             =  pe_inst[50].pe__stu__oob_data  ;

  assign   pe51__stu__valid                =  pe_inst[51].pe__stu__valid     ;
  assign   pe51__stu__cntl                 =  pe_inst[51].pe__stu__cntl      ;
  assign   pe_inst[51].stu__pe__ready      =  stu__pe51__ready               ;
  assign   pe51__stu__type                 =  pe_inst[51].pe__stu__type      ;
  assign   pe51__stu__data                 =  pe_inst[51].pe__stu__data      ;
  assign   pe51__stu__oob_data             =  pe_inst[51].pe__stu__oob_data  ;

  assign   pe52__stu__valid                =  pe_inst[52].pe__stu__valid     ;
  assign   pe52__stu__cntl                 =  pe_inst[52].pe__stu__cntl      ;
  assign   pe_inst[52].stu__pe__ready      =  stu__pe52__ready               ;
  assign   pe52__stu__type                 =  pe_inst[52].pe__stu__type      ;
  assign   pe52__stu__data                 =  pe_inst[52].pe__stu__data      ;
  assign   pe52__stu__oob_data             =  pe_inst[52].pe__stu__oob_data  ;

  assign   pe53__stu__valid                =  pe_inst[53].pe__stu__valid     ;
  assign   pe53__stu__cntl                 =  pe_inst[53].pe__stu__cntl      ;
  assign   pe_inst[53].stu__pe__ready      =  stu__pe53__ready               ;
  assign   pe53__stu__type                 =  pe_inst[53].pe__stu__type      ;
  assign   pe53__stu__data                 =  pe_inst[53].pe__stu__data      ;
  assign   pe53__stu__oob_data             =  pe_inst[53].pe__stu__oob_data  ;

  assign   pe54__stu__valid                =  pe_inst[54].pe__stu__valid     ;
  assign   pe54__stu__cntl                 =  pe_inst[54].pe__stu__cntl      ;
  assign   pe_inst[54].stu__pe__ready      =  stu__pe54__ready               ;
  assign   pe54__stu__type                 =  pe_inst[54].pe__stu__type      ;
  assign   pe54__stu__data                 =  pe_inst[54].pe__stu__data      ;
  assign   pe54__stu__oob_data             =  pe_inst[54].pe__stu__oob_data  ;

  assign   pe55__stu__valid                =  pe_inst[55].pe__stu__valid     ;
  assign   pe55__stu__cntl                 =  pe_inst[55].pe__stu__cntl      ;
  assign   pe_inst[55].stu__pe__ready      =  stu__pe55__ready               ;
  assign   pe55__stu__type                 =  pe_inst[55].pe__stu__type      ;
  assign   pe55__stu__data                 =  pe_inst[55].pe__stu__data      ;
  assign   pe55__stu__oob_data             =  pe_inst[55].pe__stu__oob_data  ;

  assign   pe56__stu__valid                =  pe_inst[56].pe__stu__valid     ;
  assign   pe56__stu__cntl                 =  pe_inst[56].pe__stu__cntl      ;
  assign   pe_inst[56].stu__pe__ready      =  stu__pe56__ready               ;
  assign   pe56__stu__type                 =  pe_inst[56].pe__stu__type      ;
  assign   pe56__stu__data                 =  pe_inst[56].pe__stu__data      ;
  assign   pe56__stu__oob_data             =  pe_inst[56].pe__stu__oob_data  ;

  assign   pe57__stu__valid                =  pe_inst[57].pe__stu__valid     ;
  assign   pe57__stu__cntl                 =  pe_inst[57].pe__stu__cntl      ;
  assign   pe_inst[57].stu__pe__ready      =  stu__pe57__ready               ;
  assign   pe57__stu__type                 =  pe_inst[57].pe__stu__type      ;
  assign   pe57__stu__data                 =  pe_inst[57].pe__stu__data      ;
  assign   pe57__stu__oob_data             =  pe_inst[57].pe__stu__oob_data  ;

  assign   pe58__stu__valid                =  pe_inst[58].pe__stu__valid     ;
  assign   pe58__stu__cntl                 =  pe_inst[58].pe__stu__cntl      ;
  assign   pe_inst[58].stu__pe__ready      =  stu__pe58__ready               ;
  assign   pe58__stu__type                 =  pe_inst[58].pe__stu__type      ;
  assign   pe58__stu__data                 =  pe_inst[58].pe__stu__data      ;
  assign   pe58__stu__oob_data             =  pe_inst[58].pe__stu__oob_data  ;

  assign   pe59__stu__valid                =  pe_inst[59].pe__stu__valid     ;
  assign   pe59__stu__cntl                 =  pe_inst[59].pe__stu__cntl      ;
  assign   pe_inst[59].stu__pe__ready      =  stu__pe59__ready               ;
  assign   pe59__stu__type                 =  pe_inst[59].pe__stu__type      ;
  assign   pe59__stu__data                 =  pe_inst[59].pe__stu__data      ;
  assign   pe59__stu__oob_data             =  pe_inst[59].pe__stu__oob_data  ;

  assign   pe60__stu__valid                =  pe_inst[60].pe__stu__valid     ;
  assign   pe60__stu__cntl                 =  pe_inst[60].pe__stu__cntl      ;
  assign   pe_inst[60].stu__pe__ready      =  stu__pe60__ready               ;
  assign   pe60__stu__type                 =  pe_inst[60].pe__stu__type      ;
  assign   pe60__stu__data                 =  pe_inst[60].pe__stu__data      ;
  assign   pe60__stu__oob_data             =  pe_inst[60].pe__stu__oob_data  ;

  assign   pe61__stu__valid                =  pe_inst[61].pe__stu__valid     ;
  assign   pe61__stu__cntl                 =  pe_inst[61].pe__stu__cntl      ;
  assign   pe_inst[61].stu__pe__ready      =  stu__pe61__ready               ;
  assign   pe61__stu__type                 =  pe_inst[61].pe__stu__type      ;
  assign   pe61__stu__data                 =  pe_inst[61].pe__stu__data      ;
  assign   pe61__stu__oob_data             =  pe_inst[61].pe__stu__oob_data  ;

  assign   pe62__stu__valid                =  pe_inst[62].pe__stu__valid     ;
  assign   pe62__stu__cntl                 =  pe_inst[62].pe__stu__cntl      ;
  assign   pe_inst[62].stu__pe__ready      =  stu__pe62__ready               ;
  assign   pe62__stu__type                 =  pe_inst[62].pe__stu__type      ;
  assign   pe62__stu__data                 =  pe_inst[62].pe__stu__data      ;
  assign   pe62__stu__oob_data             =  pe_inst[62].pe__stu__oob_data  ;

  assign   pe63__stu__valid                =  pe_inst[63].pe__stu__valid     ;
  assign   pe63__stu__cntl                 =  pe_inst[63].pe__stu__cntl      ;
  assign   pe_inst[63].stu__pe__ready      =  stu__pe63__ready               ;
  assign   pe63__stu__type                 =  pe_inst[63].pe__stu__type      ;
  assign   pe63__stu__data                 =  pe_inst[63].pe__stu__data      ;
  assign   pe63__stu__oob_data             =  pe_inst[63].pe__stu__oob_data  ;

