
`define NOC_CONT_PE0_PORT0_DESTINATION_PE_BITMASK  'b1111111011111110111111101111111011111110111111101111111011111110
`define NOC_CONT_PE0_PORT1_DESTINATION_PE_BITMASK  'b0000000100000001000000010000000100000001000000010000000100000000
`define NOC_CONT_PE0_PORT2_DESTINATION_PE_BITMASK  'd0
`define NOC_CONT_PE0_PORT3_DESTINATION_PE_BITMASK  'd0
`define NOC_CONT_PE1_PORT0_DESTINATION_PE_BITMASK  'b1111110011111100111111001111110011111100111111001111110011111100
`define NOC_CONT_PE1_PORT1_DESTINATION_PE_BITMASK  'b0000001000000010000000100000001000000010000000100000001000000000
`define NOC_CONT_PE1_PORT2_DESTINATION_PE_BITMASK  'b0000000100000001000000010000000100000001000000010000000100000001
`define NOC_CONT_PE1_PORT3_DESTINATION_PE_BITMASK  'd0
`define NOC_CONT_PE2_PORT0_DESTINATION_PE_BITMASK  'b1111100011111000111110001111100011111000111110001111100011111000
`define NOC_CONT_PE2_PORT1_DESTINATION_PE_BITMASK  'b0000010000000100000001000000010000000100000001000000010000000000
`define NOC_CONT_PE2_PORT2_DESTINATION_PE_BITMASK  'b0000001100000011000000110000001100000011000000110000001100000011
`define NOC_CONT_PE2_PORT3_DESTINATION_PE_BITMASK  'd0
`define NOC_CONT_PE3_PORT0_DESTINATION_PE_BITMASK  'b1111000011110000111100001111000011110000111100001111000011110000
`define NOC_CONT_PE3_PORT1_DESTINATION_PE_BITMASK  'b0000100000001000000010000000100000001000000010000000100000000000
`define NOC_CONT_PE3_PORT2_DESTINATION_PE_BITMASK  'b0000011100000111000001110000011100000111000001110000011100000111
`define NOC_CONT_PE3_PORT3_DESTINATION_PE_BITMASK  'd0
`define NOC_CONT_PE4_PORT0_DESTINATION_PE_BITMASK  'b1110000011100000111000001110000011100000111000001110000011100000
`define NOC_CONT_PE4_PORT1_DESTINATION_PE_BITMASK  'b0001000000010000000100000001000000010000000100000001000000000000
`define NOC_CONT_PE4_PORT2_DESTINATION_PE_BITMASK  'b0000111100001111000011110000111100001111000011110000111100001111
`define NOC_CONT_PE4_PORT3_DESTINATION_PE_BITMASK  'd0
`define NOC_CONT_PE5_PORT0_DESTINATION_PE_BITMASK  'b1100000011000000110000001100000011000000110000001100000011000000
`define NOC_CONT_PE5_PORT1_DESTINATION_PE_BITMASK  'b0010000000100000001000000010000000100000001000000010000000000000
`define NOC_CONT_PE5_PORT2_DESTINATION_PE_BITMASK  'b0001111100011111000111110001111100011111000111110001111100011111
`define NOC_CONT_PE5_PORT3_DESTINATION_PE_BITMASK  'd0
`define NOC_CONT_PE6_PORT0_DESTINATION_PE_BITMASK  'b1000000010000000100000001000000010000000100000001000000010000000
`define NOC_CONT_PE6_PORT1_DESTINATION_PE_BITMASK  'b0100000001000000010000000100000001000000010000000100000000000000
`define NOC_CONT_PE6_PORT2_DESTINATION_PE_BITMASK  'b0011111100111111001111110011111100111111001111110011111100111111
`define NOC_CONT_PE6_PORT3_DESTINATION_PE_BITMASK  'd0
`define NOC_CONT_PE7_PORT0_DESTINATION_PE_BITMASK  'b1000000010000000100000001000000010000000100000001000000000000000
`define NOC_CONT_PE7_PORT1_DESTINATION_PE_BITMASK  'b0111111101111111011111110111111101111111011111110111111101111111
`define NOC_CONT_PE7_PORT2_DESTINATION_PE_BITMASK  'd0
`define NOC_CONT_PE7_PORT3_DESTINATION_PE_BITMASK  'd0
`define NOC_CONT_PE8_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000000000000000000000000000011111111
`define NOC_CONT_PE8_PORT1_DESTINATION_PE_BITMASK  'b1111111011111110111111101111111011111110111111101111111000000000
`define NOC_CONT_PE8_PORT2_DESTINATION_PE_BITMASK  'b0000000100000001000000010000000100000001000000010000000000000000
`define NOC_CONT_PE8_PORT3_DESTINATION_PE_BITMASK  'd0
`define NOC_CONT_PE9_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000000000000000000000000000011111111
`define NOC_CONT_PE9_PORT1_DESTINATION_PE_BITMASK  'b1111110011111100111111001111110011111100111111001111110000000000
`define NOC_CONT_PE9_PORT2_DESTINATION_PE_BITMASK  'b0000001000000010000000100000001000000010000000100000000000000000
`define NOC_CONT_PE9_PORT3_DESTINATION_PE_BITMASK  'b0000000100000001000000010000000100000001000000010000000100000000
`define NOC_CONT_PE10_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000000000000000000000000000011111111
`define NOC_CONT_PE10_PORT1_DESTINATION_PE_BITMASK  'b1111100011111000111110001111100011111000111110001111100000000000
`define NOC_CONT_PE10_PORT2_DESTINATION_PE_BITMASK  'b0000010000000100000001000000010000000100000001000000000000000000
`define NOC_CONT_PE10_PORT3_DESTINATION_PE_BITMASK  'b0000001100000011000000110000001100000011000000110000001100000000
`define NOC_CONT_PE11_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000000000000000000000000000011111111
`define NOC_CONT_PE11_PORT1_DESTINATION_PE_BITMASK  'b1111000011110000111100001111000011110000111100001111000000000000
`define NOC_CONT_PE11_PORT2_DESTINATION_PE_BITMASK  'b0000100000001000000010000000100000001000000010000000000000000000
`define NOC_CONT_PE11_PORT3_DESTINATION_PE_BITMASK  'b0000011100000111000001110000011100000111000001110000011100000000
`define NOC_CONT_PE12_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000000000000000000000000000011111111
`define NOC_CONT_PE12_PORT1_DESTINATION_PE_BITMASK  'b1110000011100000111000001110000011100000111000001110000000000000
`define NOC_CONT_PE12_PORT2_DESTINATION_PE_BITMASK  'b0001000000010000000100000001000000010000000100000000000000000000
`define NOC_CONT_PE12_PORT3_DESTINATION_PE_BITMASK  'b0000111100001111000011110000111100001111000011110000111100000000
`define NOC_CONT_PE13_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000000000000000000000000000011111111
`define NOC_CONT_PE13_PORT1_DESTINATION_PE_BITMASK  'b1100000011000000110000001100000011000000110000001100000000000000
`define NOC_CONT_PE13_PORT2_DESTINATION_PE_BITMASK  'b0010000000100000001000000010000000100000001000000000000000000000
`define NOC_CONT_PE13_PORT3_DESTINATION_PE_BITMASK  'b0001111100011111000111110001111100011111000111110001111100000000
`define NOC_CONT_PE14_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000000000000000000000000000011111111
`define NOC_CONT_PE14_PORT1_DESTINATION_PE_BITMASK  'b1000000010000000100000001000000010000000100000001000000000000000
`define NOC_CONT_PE14_PORT2_DESTINATION_PE_BITMASK  'b0100000001000000010000000100000001000000010000000000000000000000
`define NOC_CONT_PE14_PORT3_DESTINATION_PE_BITMASK  'b0011111100111111001111110011111100111111001111110011111100000000
`define NOC_CONT_PE15_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000000000000000000000000000011111111
`define NOC_CONT_PE15_PORT1_DESTINATION_PE_BITMASK  'b1000000010000000100000001000000010000000100000000000000000000000
`define NOC_CONT_PE15_PORT2_DESTINATION_PE_BITMASK  'b0111111101111111011111110111111101111111011111110111111100000000
`define NOC_CONT_PE15_PORT3_DESTINATION_PE_BITMASK  'd0
`define NOC_CONT_PE16_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000000000000000000001111111111111111
`define NOC_CONT_PE16_PORT1_DESTINATION_PE_BITMASK  'b1111111011111110111111101111111011111110111111100000000000000000
`define NOC_CONT_PE16_PORT2_DESTINATION_PE_BITMASK  'b0000000100000001000000010000000100000001000000000000000000000000
`define NOC_CONT_PE16_PORT3_DESTINATION_PE_BITMASK  'd0
`define NOC_CONT_PE17_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000000000000000000001111111111111111
`define NOC_CONT_PE17_PORT1_DESTINATION_PE_BITMASK  'b1111110011111100111111001111110011111100111111000000000000000000
`define NOC_CONT_PE17_PORT2_DESTINATION_PE_BITMASK  'b0000001000000010000000100000001000000010000000000000000000000000
`define NOC_CONT_PE17_PORT3_DESTINATION_PE_BITMASK  'b0000000100000001000000010000000100000001000000010000000000000000
`define NOC_CONT_PE18_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000000000000000000001111111111111111
`define NOC_CONT_PE18_PORT1_DESTINATION_PE_BITMASK  'b1111100011111000111110001111100011111000111110000000000000000000
`define NOC_CONT_PE18_PORT2_DESTINATION_PE_BITMASK  'b0000010000000100000001000000010000000100000000000000000000000000
`define NOC_CONT_PE18_PORT3_DESTINATION_PE_BITMASK  'b0000001100000011000000110000001100000011000000110000000000000000
`define NOC_CONT_PE19_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000000000000000000001111111111111111
`define NOC_CONT_PE19_PORT1_DESTINATION_PE_BITMASK  'b1111000011110000111100001111000011110000111100000000000000000000
`define NOC_CONT_PE19_PORT2_DESTINATION_PE_BITMASK  'b0000100000001000000010000000100000001000000000000000000000000000
`define NOC_CONT_PE19_PORT3_DESTINATION_PE_BITMASK  'b0000011100000111000001110000011100000111000001110000000000000000
`define NOC_CONT_PE20_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000000000000000000001111111111111111
`define NOC_CONT_PE20_PORT1_DESTINATION_PE_BITMASK  'b1110000011100000111000001110000011100000111000000000000000000000
`define NOC_CONT_PE20_PORT2_DESTINATION_PE_BITMASK  'b0001000000010000000100000001000000010000000000000000000000000000
`define NOC_CONT_PE20_PORT3_DESTINATION_PE_BITMASK  'b0000111100001111000011110000111100001111000011110000000000000000
`define NOC_CONT_PE21_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000000000000000000001111111111111111
`define NOC_CONT_PE21_PORT1_DESTINATION_PE_BITMASK  'b1100000011000000110000001100000011000000110000000000000000000000
`define NOC_CONT_PE21_PORT2_DESTINATION_PE_BITMASK  'b0010000000100000001000000010000000100000000000000000000000000000
`define NOC_CONT_PE21_PORT3_DESTINATION_PE_BITMASK  'b0001111100011111000111110001111100011111000111110000000000000000
`define NOC_CONT_PE22_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000000000000000000001111111111111111
`define NOC_CONT_PE22_PORT1_DESTINATION_PE_BITMASK  'b1000000010000000100000001000000010000000100000000000000000000000
`define NOC_CONT_PE22_PORT2_DESTINATION_PE_BITMASK  'b0100000001000000010000000100000001000000000000000000000000000000
`define NOC_CONT_PE22_PORT3_DESTINATION_PE_BITMASK  'b0011111100111111001111110011111100111111001111110000000000000000
`define NOC_CONT_PE23_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000000000000000000001111111111111111
`define NOC_CONT_PE23_PORT1_DESTINATION_PE_BITMASK  'b1000000010000000100000001000000010000000000000000000000000000000
`define NOC_CONT_PE23_PORT2_DESTINATION_PE_BITMASK  'b0111111101111111011111110111111101111111011111110000000000000000
`define NOC_CONT_PE23_PORT3_DESTINATION_PE_BITMASK  'd0
`define NOC_CONT_PE24_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000000000000111111111111111111111111
`define NOC_CONT_PE24_PORT1_DESTINATION_PE_BITMASK  'b1111111011111110111111101111111011111110000000000000000000000000
`define NOC_CONT_PE24_PORT2_DESTINATION_PE_BITMASK  'b0000000100000001000000010000000100000000000000000000000000000000
`define NOC_CONT_PE24_PORT3_DESTINATION_PE_BITMASK  'd0
`define NOC_CONT_PE25_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000000000000111111111111111111111111
`define NOC_CONT_PE25_PORT1_DESTINATION_PE_BITMASK  'b1111110011111100111111001111110011111100000000000000000000000000
`define NOC_CONT_PE25_PORT2_DESTINATION_PE_BITMASK  'b0000001000000010000000100000001000000000000000000000000000000000
`define NOC_CONT_PE25_PORT3_DESTINATION_PE_BITMASK  'b0000000100000001000000010000000100000001000000000000000000000000
`define NOC_CONT_PE26_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000000000000111111111111111111111111
`define NOC_CONT_PE26_PORT1_DESTINATION_PE_BITMASK  'b1111100011111000111110001111100011111000000000000000000000000000
`define NOC_CONT_PE26_PORT2_DESTINATION_PE_BITMASK  'b0000010000000100000001000000010000000000000000000000000000000000
`define NOC_CONT_PE26_PORT3_DESTINATION_PE_BITMASK  'b0000001100000011000000110000001100000011000000000000000000000000
`define NOC_CONT_PE27_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000000000000111111111111111111111111
`define NOC_CONT_PE27_PORT1_DESTINATION_PE_BITMASK  'b1111000011110000111100001111000011110000000000000000000000000000
`define NOC_CONT_PE27_PORT2_DESTINATION_PE_BITMASK  'b0000100000001000000010000000100000000000000000000000000000000000
`define NOC_CONT_PE27_PORT3_DESTINATION_PE_BITMASK  'b0000011100000111000001110000011100000111000000000000000000000000
`define NOC_CONT_PE28_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000000000000111111111111111111111111
`define NOC_CONT_PE28_PORT1_DESTINATION_PE_BITMASK  'b1110000011100000111000001110000011100000000000000000000000000000
`define NOC_CONT_PE28_PORT2_DESTINATION_PE_BITMASK  'b0001000000010000000100000001000000000000000000000000000000000000
`define NOC_CONT_PE28_PORT3_DESTINATION_PE_BITMASK  'b0000111100001111000011110000111100001111000000000000000000000000
`define NOC_CONT_PE29_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000000000000111111111111111111111111
`define NOC_CONT_PE29_PORT1_DESTINATION_PE_BITMASK  'b1100000011000000110000001100000011000000000000000000000000000000
`define NOC_CONT_PE29_PORT2_DESTINATION_PE_BITMASK  'b0010000000100000001000000010000000000000000000000000000000000000
`define NOC_CONT_PE29_PORT3_DESTINATION_PE_BITMASK  'b0001111100011111000111110001111100011111000000000000000000000000
`define NOC_CONT_PE30_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000000000000111111111111111111111111
`define NOC_CONT_PE30_PORT1_DESTINATION_PE_BITMASK  'b1000000010000000100000001000000010000000000000000000000000000000
`define NOC_CONT_PE30_PORT2_DESTINATION_PE_BITMASK  'b0100000001000000010000000100000000000000000000000000000000000000
`define NOC_CONT_PE30_PORT3_DESTINATION_PE_BITMASK  'b0011111100111111001111110011111100111111000000000000000000000000
`define NOC_CONT_PE31_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000000000000111111111111111111111111
`define NOC_CONT_PE31_PORT1_DESTINATION_PE_BITMASK  'b1000000010000000100000001000000000000000000000000000000000000000
`define NOC_CONT_PE31_PORT2_DESTINATION_PE_BITMASK  'b0111111101111111011111110111111101111111000000000000000000000000
`define NOC_CONT_PE31_PORT3_DESTINATION_PE_BITMASK  'd0
`define NOC_CONT_PE32_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000011111111111111111111111111111111
`define NOC_CONT_PE32_PORT1_DESTINATION_PE_BITMASK  'b1111111011111110111111101111111000000000000000000000000000000000
`define NOC_CONT_PE32_PORT2_DESTINATION_PE_BITMASK  'b0000000100000001000000010000000000000000000000000000000000000000
`define NOC_CONT_PE32_PORT3_DESTINATION_PE_BITMASK  'd0
`define NOC_CONT_PE33_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000011111111111111111111111111111111
`define NOC_CONT_PE33_PORT1_DESTINATION_PE_BITMASK  'b1111110011111100111111001111110000000000000000000000000000000000
`define NOC_CONT_PE33_PORT2_DESTINATION_PE_BITMASK  'b0000001000000010000000100000000000000000000000000000000000000000
`define NOC_CONT_PE33_PORT3_DESTINATION_PE_BITMASK  'b0000000100000001000000010000000100000000000000000000000000000000
`define NOC_CONT_PE34_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000011111111111111111111111111111111
`define NOC_CONT_PE34_PORT1_DESTINATION_PE_BITMASK  'b1111100011111000111110001111100000000000000000000000000000000000
`define NOC_CONT_PE34_PORT2_DESTINATION_PE_BITMASK  'b0000010000000100000001000000000000000000000000000000000000000000
`define NOC_CONT_PE34_PORT3_DESTINATION_PE_BITMASK  'b0000001100000011000000110000001100000000000000000000000000000000
`define NOC_CONT_PE35_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000011111111111111111111111111111111
`define NOC_CONT_PE35_PORT1_DESTINATION_PE_BITMASK  'b1111000011110000111100001111000000000000000000000000000000000000
`define NOC_CONT_PE35_PORT2_DESTINATION_PE_BITMASK  'b0000100000001000000010000000000000000000000000000000000000000000
`define NOC_CONT_PE35_PORT3_DESTINATION_PE_BITMASK  'b0000011100000111000001110000011100000000000000000000000000000000
`define NOC_CONT_PE36_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000011111111111111111111111111111111
`define NOC_CONT_PE36_PORT1_DESTINATION_PE_BITMASK  'b1110000011100000111000001110000000000000000000000000000000000000
`define NOC_CONT_PE36_PORT2_DESTINATION_PE_BITMASK  'b0001000000010000000100000000000000000000000000000000000000000000
`define NOC_CONT_PE36_PORT3_DESTINATION_PE_BITMASK  'b0000111100001111000011110000111100000000000000000000000000000000
`define NOC_CONT_PE37_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000011111111111111111111111111111111
`define NOC_CONT_PE37_PORT1_DESTINATION_PE_BITMASK  'b1100000011000000110000001100000000000000000000000000000000000000
`define NOC_CONT_PE37_PORT2_DESTINATION_PE_BITMASK  'b0010000000100000001000000000000000000000000000000000000000000000
`define NOC_CONT_PE37_PORT3_DESTINATION_PE_BITMASK  'b0001111100011111000111110001111100000000000000000000000000000000
`define NOC_CONT_PE38_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000011111111111111111111111111111111
`define NOC_CONT_PE38_PORT1_DESTINATION_PE_BITMASK  'b1000000010000000100000001000000000000000000000000000000000000000
`define NOC_CONT_PE38_PORT2_DESTINATION_PE_BITMASK  'b0100000001000000010000000000000000000000000000000000000000000000
`define NOC_CONT_PE38_PORT3_DESTINATION_PE_BITMASK  'b0011111100111111001111110011111100000000000000000000000000000000
`define NOC_CONT_PE39_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000000000000011111111111111111111111111111111
`define NOC_CONT_PE39_PORT1_DESTINATION_PE_BITMASK  'b1000000010000000100000000000000000000000000000000000000000000000
`define NOC_CONT_PE39_PORT2_DESTINATION_PE_BITMASK  'b0111111101111111011111110111111100000000000000000000000000000000
`define NOC_CONT_PE39_PORT3_DESTINATION_PE_BITMASK  'd0
`define NOC_CONT_PE40_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000001111111111111111111111111111111111111111
`define NOC_CONT_PE40_PORT1_DESTINATION_PE_BITMASK  'b1111111011111110111111100000000000000000000000000000000000000000
`define NOC_CONT_PE40_PORT2_DESTINATION_PE_BITMASK  'b0000000100000001000000000000000000000000000000000000000000000000
`define NOC_CONT_PE40_PORT3_DESTINATION_PE_BITMASK  'd0
`define NOC_CONT_PE41_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000001111111111111111111111111111111111111111
`define NOC_CONT_PE41_PORT1_DESTINATION_PE_BITMASK  'b1111110011111100111111000000000000000000000000000000000000000000
`define NOC_CONT_PE41_PORT2_DESTINATION_PE_BITMASK  'b0000001000000010000000000000000000000000000000000000000000000000
`define NOC_CONT_PE41_PORT3_DESTINATION_PE_BITMASK  'b0000000100000001000000010000000000000000000000000000000000000000
`define NOC_CONT_PE42_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000001111111111111111111111111111111111111111
`define NOC_CONT_PE42_PORT1_DESTINATION_PE_BITMASK  'b1111100011111000111110000000000000000000000000000000000000000000
`define NOC_CONT_PE42_PORT2_DESTINATION_PE_BITMASK  'b0000010000000100000000000000000000000000000000000000000000000000
`define NOC_CONT_PE42_PORT3_DESTINATION_PE_BITMASK  'b0000001100000011000000110000000000000000000000000000000000000000
`define NOC_CONT_PE43_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000001111111111111111111111111111111111111111
`define NOC_CONT_PE43_PORT1_DESTINATION_PE_BITMASK  'b1111000011110000111100000000000000000000000000000000000000000000
`define NOC_CONT_PE43_PORT2_DESTINATION_PE_BITMASK  'b0000100000001000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE43_PORT3_DESTINATION_PE_BITMASK  'b0000011100000111000001110000000000000000000000000000000000000000
`define NOC_CONT_PE44_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000001111111111111111111111111111111111111111
`define NOC_CONT_PE44_PORT1_DESTINATION_PE_BITMASK  'b1110000011100000111000000000000000000000000000000000000000000000
`define NOC_CONT_PE44_PORT2_DESTINATION_PE_BITMASK  'b0001000000010000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE44_PORT3_DESTINATION_PE_BITMASK  'b0000111100001111000011110000000000000000000000000000000000000000
`define NOC_CONT_PE45_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000001111111111111111111111111111111111111111
`define NOC_CONT_PE45_PORT1_DESTINATION_PE_BITMASK  'b1100000011000000110000000000000000000000000000000000000000000000
`define NOC_CONT_PE45_PORT2_DESTINATION_PE_BITMASK  'b0010000000100000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE45_PORT3_DESTINATION_PE_BITMASK  'b0001111100011111000111110000000000000000000000000000000000000000
`define NOC_CONT_PE46_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000001111111111111111111111111111111111111111
`define NOC_CONT_PE46_PORT1_DESTINATION_PE_BITMASK  'b1000000010000000100000000000000000000000000000000000000000000000
`define NOC_CONT_PE46_PORT2_DESTINATION_PE_BITMASK  'b0100000001000000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE46_PORT3_DESTINATION_PE_BITMASK  'b0011111100111111001111110000000000000000000000000000000000000000
`define NOC_CONT_PE47_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000000000001111111111111111111111111111111111111111
`define NOC_CONT_PE47_PORT1_DESTINATION_PE_BITMASK  'b1000000010000000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE47_PORT2_DESTINATION_PE_BITMASK  'b0111111101111111011111110000000000000000000000000000000000000000
`define NOC_CONT_PE47_PORT3_DESTINATION_PE_BITMASK  'd0
`define NOC_CONT_PE48_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000111111111111111111111111111111111111111111111111
`define NOC_CONT_PE48_PORT1_DESTINATION_PE_BITMASK  'b1111111011111110000000000000000000000000000000000000000000000000
`define NOC_CONT_PE48_PORT2_DESTINATION_PE_BITMASK  'b0000000100000000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE48_PORT3_DESTINATION_PE_BITMASK  'd0
`define NOC_CONT_PE49_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000111111111111111111111111111111111111111111111111
`define NOC_CONT_PE49_PORT1_DESTINATION_PE_BITMASK  'b1111110011111100000000000000000000000000000000000000000000000000
`define NOC_CONT_PE49_PORT2_DESTINATION_PE_BITMASK  'b0000001000000000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE49_PORT3_DESTINATION_PE_BITMASK  'b0000000100000001000000000000000000000000000000000000000000000000
`define NOC_CONT_PE50_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000111111111111111111111111111111111111111111111111
`define NOC_CONT_PE50_PORT1_DESTINATION_PE_BITMASK  'b1111100011111000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE50_PORT2_DESTINATION_PE_BITMASK  'b0000010000000000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE50_PORT3_DESTINATION_PE_BITMASK  'b0000001100000011000000000000000000000000000000000000000000000000
`define NOC_CONT_PE51_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000111111111111111111111111111111111111111111111111
`define NOC_CONT_PE51_PORT1_DESTINATION_PE_BITMASK  'b1111000011110000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE51_PORT2_DESTINATION_PE_BITMASK  'b0000100000000000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE51_PORT3_DESTINATION_PE_BITMASK  'b0000011100000111000000000000000000000000000000000000000000000000
`define NOC_CONT_PE52_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000111111111111111111111111111111111111111111111111
`define NOC_CONT_PE52_PORT1_DESTINATION_PE_BITMASK  'b1110000011100000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE52_PORT2_DESTINATION_PE_BITMASK  'b0001000000000000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE52_PORT3_DESTINATION_PE_BITMASK  'b0000111100001111000000000000000000000000000000000000000000000000
`define NOC_CONT_PE53_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000111111111111111111111111111111111111111111111111
`define NOC_CONT_PE53_PORT1_DESTINATION_PE_BITMASK  'b1100000011000000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE53_PORT2_DESTINATION_PE_BITMASK  'b0010000000000000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE53_PORT3_DESTINATION_PE_BITMASK  'b0001111100011111000000000000000000000000000000000000000000000000
`define NOC_CONT_PE54_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000111111111111111111111111111111111111111111111111
`define NOC_CONT_PE54_PORT1_DESTINATION_PE_BITMASK  'b1000000010000000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE54_PORT2_DESTINATION_PE_BITMASK  'b0100000000000000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE54_PORT3_DESTINATION_PE_BITMASK  'b0011111100111111000000000000000000000000000000000000000000000000
`define NOC_CONT_PE55_PORT0_DESTINATION_PE_BITMASK  'b0000000000000000111111111111111111111111111111111111111111111111
`define NOC_CONT_PE55_PORT1_DESTINATION_PE_BITMASK  'b1000000000000000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE55_PORT2_DESTINATION_PE_BITMASK  'b0111111101111111000000000000000000000000000000000000000000000000
`define NOC_CONT_PE55_PORT3_DESTINATION_PE_BITMASK  'd0
`define NOC_CONT_PE56_PORT0_DESTINATION_PE_BITMASK  'b0000000011111111111111111111111111111111111111111111111111111111
`define NOC_CONT_PE56_PORT1_DESTINATION_PE_BITMASK  'b1111111000000000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE56_PORT2_DESTINATION_PE_BITMASK  'd0
`define NOC_CONT_PE56_PORT3_DESTINATION_PE_BITMASK  'd0
`define NOC_CONT_PE57_PORT0_DESTINATION_PE_BITMASK  'b0000000011111111111111111111111111111111111111111111111111111111
`define NOC_CONT_PE57_PORT1_DESTINATION_PE_BITMASK  'b1111110000000000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE57_PORT2_DESTINATION_PE_BITMASK  'b0000000100000000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE57_PORT3_DESTINATION_PE_BITMASK  'd0
`define NOC_CONT_PE58_PORT0_DESTINATION_PE_BITMASK  'b0000000011111111111111111111111111111111111111111111111111111111
`define NOC_CONT_PE58_PORT1_DESTINATION_PE_BITMASK  'b1111100000000000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE58_PORT2_DESTINATION_PE_BITMASK  'b0000001100000000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE58_PORT3_DESTINATION_PE_BITMASK  'd0
`define NOC_CONT_PE59_PORT0_DESTINATION_PE_BITMASK  'b0000000011111111111111111111111111111111111111111111111111111111
`define NOC_CONT_PE59_PORT1_DESTINATION_PE_BITMASK  'b1111000000000000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE59_PORT2_DESTINATION_PE_BITMASK  'b0000011100000000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE59_PORT3_DESTINATION_PE_BITMASK  'd0
`define NOC_CONT_PE60_PORT0_DESTINATION_PE_BITMASK  'b0000000011111111111111111111111111111111111111111111111111111111
`define NOC_CONT_PE60_PORT1_DESTINATION_PE_BITMASK  'b1110000000000000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE60_PORT2_DESTINATION_PE_BITMASK  'b0000111100000000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE60_PORT3_DESTINATION_PE_BITMASK  'd0
`define NOC_CONT_PE61_PORT0_DESTINATION_PE_BITMASK  'b0000000011111111111111111111111111111111111111111111111111111111
`define NOC_CONT_PE61_PORT1_DESTINATION_PE_BITMASK  'b1100000000000000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE61_PORT2_DESTINATION_PE_BITMASK  'b0001111100000000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE61_PORT3_DESTINATION_PE_BITMASK  'd0
`define NOC_CONT_PE62_PORT0_DESTINATION_PE_BITMASK  'b0000000011111111111111111111111111111111111111111111111111111111
`define NOC_CONT_PE62_PORT1_DESTINATION_PE_BITMASK  'b1000000000000000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE62_PORT2_DESTINATION_PE_BITMASK  'b0011111100000000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE62_PORT3_DESTINATION_PE_BITMASK  'd0
`define NOC_CONT_PE63_PORT0_DESTINATION_PE_BITMASK  'b0000000011111111111111111111111111111111111111111111111111111111
`define NOC_CONT_PE63_PORT1_DESTINATION_PE_BITMASK  'b0111111100000000000000000000000000000000000000000000000000000000
`define NOC_CONT_PE63_PORT2_DESTINATION_PE_BITMASK  'd0
`define NOC_CONT_PE63_PORT3_DESTINATION_PE_BITMASK  'd0
