
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr0__std__oob_cntl            ;
  output                                          mgr0__std__oob_valid           ;
  input                                           std__mgr0__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr0__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr0__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr1__std__oob_cntl            ;
  output                                          mgr1__std__oob_valid           ;
  input                                           std__mgr1__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr1__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr1__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr2__std__oob_cntl            ;
  output                                          mgr2__std__oob_valid           ;
  input                                           std__mgr2__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr2__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr2__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr3__std__oob_cntl            ;
  output                                          mgr3__std__oob_valid           ;
  input                                           std__mgr3__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr3__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr3__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr4__std__oob_cntl            ;
  output                                          mgr4__std__oob_valid           ;
  input                                           std__mgr4__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr4__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr4__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr5__std__oob_cntl            ;
  output                                          mgr5__std__oob_valid           ;
  input                                           std__mgr5__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr5__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr5__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr6__std__oob_cntl            ;
  output                                          mgr6__std__oob_valid           ;
  input                                           std__mgr6__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr6__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr6__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr7__std__oob_cntl            ;
  output                                          mgr7__std__oob_valid           ;
  input                                           std__mgr7__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr7__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr7__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr8__std__oob_cntl            ;
  output                                          mgr8__std__oob_valid           ;
  input                                           std__mgr8__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr8__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr8__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr9__std__oob_cntl            ;
  output                                          mgr9__std__oob_valid           ;
  input                                           std__mgr9__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr9__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr9__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr10__std__oob_cntl            ;
  output                                          mgr10__std__oob_valid           ;
  input                                           std__mgr10__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr10__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr10__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr11__std__oob_cntl            ;
  output                                          mgr11__std__oob_valid           ;
  input                                           std__mgr11__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr11__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr11__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr12__std__oob_cntl            ;
  output                                          mgr12__std__oob_valid           ;
  input                                           std__mgr12__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr12__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr12__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr13__std__oob_cntl            ;
  output                                          mgr13__std__oob_valid           ;
  input                                           std__mgr13__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr13__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr13__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr14__std__oob_cntl            ;
  output                                          mgr14__std__oob_valid           ;
  input                                           std__mgr14__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr14__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr14__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr15__std__oob_cntl            ;
  output                                          mgr15__std__oob_valid           ;
  input                                           std__mgr15__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr15__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr15__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr16__std__oob_cntl            ;
  output                                          mgr16__std__oob_valid           ;
  input                                           std__mgr16__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr16__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr16__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr17__std__oob_cntl            ;
  output                                          mgr17__std__oob_valid           ;
  input                                           std__mgr17__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr17__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr17__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr18__std__oob_cntl            ;
  output                                          mgr18__std__oob_valid           ;
  input                                           std__mgr18__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr18__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr18__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr19__std__oob_cntl            ;
  output                                          mgr19__std__oob_valid           ;
  input                                           std__mgr19__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr19__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr19__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr20__std__oob_cntl            ;
  output                                          mgr20__std__oob_valid           ;
  input                                           std__mgr20__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr20__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr20__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr21__std__oob_cntl            ;
  output                                          mgr21__std__oob_valid           ;
  input                                           std__mgr21__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr21__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr21__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr22__std__oob_cntl            ;
  output                                          mgr22__std__oob_valid           ;
  input                                           std__mgr22__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr22__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr22__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr23__std__oob_cntl            ;
  output                                          mgr23__std__oob_valid           ;
  input                                           std__mgr23__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr23__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr23__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr24__std__oob_cntl            ;
  output                                          mgr24__std__oob_valid           ;
  input                                           std__mgr24__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr24__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr24__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr25__std__oob_cntl            ;
  output                                          mgr25__std__oob_valid           ;
  input                                           std__mgr25__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr25__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr25__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr26__std__oob_cntl            ;
  output                                          mgr26__std__oob_valid           ;
  input                                           std__mgr26__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr26__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr26__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr27__std__oob_cntl            ;
  output                                          mgr27__std__oob_valid           ;
  input                                           std__mgr27__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr27__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr27__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr28__std__oob_cntl            ;
  output                                          mgr28__std__oob_valid           ;
  input                                           std__mgr28__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr28__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr28__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr29__std__oob_cntl            ;
  output                                          mgr29__std__oob_valid           ;
  input                                           std__mgr29__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr29__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr29__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr30__std__oob_cntl            ;
  output                                          mgr30__std__oob_valid           ;
  input                                           std__mgr30__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr30__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr30__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr31__std__oob_cntl            ;
  output                                          mgr31__std__oob_valid           ;
  input                                           std__mgr31__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr31__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr31__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr32__std__oob_cntl            ;
  output                                          mgr32__std__oob_valid           ;
  input                                           std__mgr32__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr32__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr32__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr33__std__oob_cntl            ;
  output                                          mgr33__std__oob_valid           ;
  input                                           std__mgr33__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr33__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr33__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr34__std__oob_cntl            ;
  output                                          mgr34__std__oob_valid           ;
  input                                           std__mgr34__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr34__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr34__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr35__std__oob_cntl            ;
  output                                          mgr35__std__oob_valid           ;
  input                                           std__mgr35__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr35__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr35__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr36__std__oob_cntl            ;
  output                                          mgr36__std__oob_valid           ;
  input                                           std__mgr36__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr36__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr36__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr37__std__oob_cntl            ;
  output                                          mgr37__std__oob_valid           ;
  input                                           std__mgr37__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr37__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr37__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr38__std__oob_cntl            ;
  output                                          mgr38__std__oob_valid           ;
  input                                           std__mgr38__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr38__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr38__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr39__std__oob_cntl            ;
  output                                          mgr39__std__oob_valid           ;
  input                                           std__mgr39__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr39__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr39__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr40__std__oob_cntl            ;
  output                                          mgr40__std__oob_valid           ;
  input                                           std__mgr40__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr40__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr40__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr41__std__oob_cntl            ;
  output                                          mgr41__std__oob_valid           ;
  input                                           std__mgr41__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr41__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr41__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr42__std__oob_cntl            ;
  output                                          mgr42__std__oob_valid           ;
  input                                           std__mgr42__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr42__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr42__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr43__std__oob_cntl            ;
  output                                          mgr43__std__oob_valid           ;
  input                                           std__mgr43__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr43__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr43__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr44__std__oob_cntl            ;
  output                                          mgr44__std__oob_valid           ;
  input                                           std__mgr44__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr44__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr44__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr45__std__oob_cntl            ;
  output                                          mgr45__std__oob_valid           ;
  input                                           std__mgr45__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr45__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr45__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr46__std__oob_cntl            ;
  output                                          mgr46__std__oob_valid           ;
  input                                           std__mgr46__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr46__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr46__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr47__std__oob_cntl            ;
  output                                          mgr47__std__oob_valid           ;
  input                                           std__mgr47__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr47__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr47__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr48__std__oob_cntl            ;
  output                                          mgr48__std__oob_valid           ;
  input                                           std__mgr48__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr48__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr48__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr49__std__oob_cntl            ;
  output                                          mgr49__std__oob_valid           ;
  input                                           std__mgr49__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr49__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr49__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr50__std__oob_cntl            ;
  output                                          mgr50__std__oob_valid           ;
  input                                           std__mgr50__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr50__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr50__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr51__std__oob_cntl            ;
  output                                          mgr51__std__oob_valid           ;
  input                                           std__mgr51__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr51__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr51__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr52__std__oob_cntl            ;
  output                                          mgr52__std__oob_valid           ;
  input                                           std__mgr52__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr52__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr52__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr53__std__oob_cntl            ;
  output                                          mgr53__std__oob_valid           ;
  input                                           std__mgr53__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr53__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr53__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr54__std__oob_cntl            ;
  output                                          mgr54__std__oob_valid           ;
  input                                           std__mgr54__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr54__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr54__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr55__std__oob_cntl            ;
  output                                          mgr55__std__oob_valid           ;
  input                                           std__mgr55__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr55__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr55__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr56__std__oob_cntl            ;
  output                                          mgr56__std__oob_valid           ;
  input                                           std__mgr56__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr56__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr56__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr57__std__oob_cntl            ;
  output                                          mgr57__std__oob_valid           ;
  input                                           std__mgr57__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr57__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr57__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr58__std__oob_cntl            ;
  output                                          mgr58__std__oob_valid           ;
  input                                           std__mgr58__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr58__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr58__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr59__std__oob_cntl            ;
  output                                          mgr59__std__oob_valid           ;
  input                                           std__mgr59__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr59__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr59__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr60__std__oob_cntl            ;
  output                                          mgr60__std__oob_valid           ;
  input                                           std__mgr60__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr60__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr60__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr61__std__oob_cntl            ;
  output                                          mgr61__std__oob_valid           ;
  input                                           std__mgr61__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr61__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr61__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr62__std__oob_cntl            ;
  output                                          mgr62__std__oob_valid           ;
  input                                           std__mgr62__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr62__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr62__std__oob_data            ;
  // OOB controls how the lanes are interpreted                                  
  output  [`COMMON_STD_INTF_CNTL_RANGE     ]      mgr63__std__oob_cntl            ;
  output                                          mgr63__std__oob_valid           ;
  input                                           std__mgr63__oob_ready           ;
  output  [`STACK_DOWN_OOB_INTF_TYPE_RANGE ]      mgr63__std__oob_type            ;
  output  [`STACK_DOWN_OOB_INTF_DATA_RANGE ]      mgr63__std__oob_data            ;