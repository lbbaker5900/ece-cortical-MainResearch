
    0 :
      begin
        to_Stu_Fifo[0].write_data   <= {simd__sui__regs[3],  
                                        simd__sui__regs[2],  
                                        simd__sui__regs[1],  
                                        simd__sui__regs[0]}; 
      end 
    1 :
      begin
        to_Stu_Fifo[0].write_data   <= {simd__sui__regs[7],  
                                        simd__sui__regs[6],  
                                        simd__sui__regs[5],  
                                        simd__sui__regs[4]}; 
      end 
    2 :
      begin
        to_Stu_Fifo[0].write_data   <= {simd__sui__regs[11],  
                                        simd__sui__regs[10],  
                                        simd__sui__regs[9],  
                                        simd__sui__regs[8]}; 
      end 
    3 :
      begin
        to_Stu_Fifo[0].write_data   <= {simd__sui__regs[15],  
                                        simd__sui__regs[14],  
                                        simd__sui__regs[13],  
                                        simd__sui__regs[12]}; 
      end 
    4 :
      begin
        to_Stu_Fifo[0].write_data   <= {simd__sui__regs[19],  
                                        simd__sui__regs[18],  
                                        simd__sui__regs[17],  
                                        simd__sui__regs[16]}; 
      end 
    5 :
      begin
        to_Stu_Fifo[0].write_data   <= {simd__sui__regs[23],  
                                        simd__sui__regs[22],  
                                        simd__sui__regs[21],  
                                        simd__sui__regs[20]}; 
      end 
    6 :
      begin
        to_Stu_Fifo[0].write_data   <= {simd__sui__regs[27],  
                                        simd__sui__regs[26],  
                                        simd__sui__regs[25],  
                                        simd__sui__regs[24]}; 
      end 
    7 :
      begin
        to_Stu_Fifo[0].write_data   <= {simd__sui__regs[31],  
                                        simd__sui__regs[30],  
                                        simd__sui__regs[29],  
                                        simd__sui__regs[28]}; 
      end 