
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  rs0  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  rs1  ;

// Lane 0                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane0_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane0_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane0_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane0_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane0_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane0_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane0_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane0_r135  ;

// Lane 1                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane1_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane1_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane1_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane1_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane1_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane1_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane1_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane1_r135  ;

// Lane 2                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane2_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane2_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane2_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane2_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane2_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane2_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane2_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane2_r135  ;

// Lane 3                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane3_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane3_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane3_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane3_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane3_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane3_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane3_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane3_r135  ;

// Lane 4                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane4_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane4_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane4_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane4_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane4_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane4_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane4_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane4_r135  ;

// Lane 5                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane5_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane5_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane5_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane5_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane5_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane5_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane5_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane5_r135  ;

// Lane 6                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane6_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane6_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane6_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane6_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane6_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane6_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane6_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane6_r135  ;

// Lane 7                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane7_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane7_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane7_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane7_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane7_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane7_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane7_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane7_r135  ;

// Lane 8                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane8_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane8_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane8_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane8_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane8_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane8_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane8_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane8_r135  ;

// Lane 9                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane9_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane9_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane9_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane9_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane9_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane9_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane9_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane9_r135  ;

// Lane 10                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane10_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane10_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane10_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane10_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane10_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane10_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane10_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane10_r135  ;

// Lane 11                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane11_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane11_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane11_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane11_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane11_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane11_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane11_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane11_r135  ;

// Lane 12                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane12_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane12_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane12_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane12_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane12_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane12_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane12_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane12_r135  ;

// Lane 13                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane13_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane13_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane13_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane13_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane13_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane13_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane13_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane13_r135  ;

// Lane 14                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane14_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane14_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane14_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane14_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane14_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane14_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane14_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane14_r135  ;

// Lane 15                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane15_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane15_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane15_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane15_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane15_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane15_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane15_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane15_r135  ;

// Lane 16                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane16_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane16_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane16_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane16_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane16_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane16_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane16_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane16_r135  ;

// Lane 17                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane17_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane17_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane17_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane17_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane17_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane17_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane17_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane17_r135  ;

// Lane 18                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane18_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane18_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane18_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane18_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane18_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane18_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane18_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane18_r135  ;

// Lane 19                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane19_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane19_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane19_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane19_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane19_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane19_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane19_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane19_r135  ;

// Lane 20                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane20_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane20_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane20_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane20_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane20_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane20_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane20_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane20_r135  ;

// Lane 21                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane21_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane21_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane21_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane21_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane21_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane21_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane21_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane21_r135  ;

// Lane 22                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane22_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane22_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane22_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane22_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane22_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane22_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane22_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane22_r135  ;

// Lane 23                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane23_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane23_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane23_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane23_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane23_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane23_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane23_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane23_r135  ;

// Lane 24                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane24_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane24_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane24_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane24_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane24_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane24_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane24_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane24_r135  ;

// Lane 25                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane25_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane25_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane25_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane25_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane25_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane25_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane25_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane25_r135  ;

// Lane 26                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane26_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane26_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane26_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane26_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane26_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane26_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane26_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane26_r135  ;

// Lane 27                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane27_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane27_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane27_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane27_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane27_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane27_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane27_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane27_r135  ;

// Lane 28                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane28_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane28_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane28_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane28_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane28_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane28_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane28_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane28_r135  ;

// Lane 29                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane29_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane29_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane29_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane29_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane29_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane29_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane29_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane29_r135  ;

// Lane 30                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane30_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane30_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane30_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane30_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane30_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane30_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane30_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane30_r135  ;

// Lane 31                 
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane31_r128  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane31_r129  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane31_r130  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane31_r131  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane31_r132  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane31_r133  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane31_r134  ;
  wire [`PE_EXEC_LANE_WIDTH_RANGE]  lane31_r135  ;
