

            // ##################################################
            // DMA Stream start addresses

            // Stream 0 start address
            force pe_array_inst.pe_inst[0].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[0].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[0].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[0].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[0].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[0].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[0].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[0].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[0].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[0].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[0].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[0].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[0].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[0].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[0].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[0].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[0].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[0].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[0].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[0].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[0].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[0].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[0].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[0].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[0].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[0].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[0].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[0].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[0].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[0].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[0].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[0].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[0].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[0].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[0].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[0].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[0].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[0].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[0].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[0].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[0].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[0].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[0].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[0].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[0].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[0].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[0].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[0].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[0].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[0].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[0].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[0].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[0].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[0].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[0].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[0].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[0].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[0].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[0].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[0].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[0].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[0].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[0].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[0].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[1].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[1].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[1].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[1].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[1].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[1].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[1].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[1].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[1].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[1].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[1].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[1].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[1].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[1].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[1].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[1].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[1].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[1].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[1].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[1].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[1].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[1].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[1].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[1].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[1].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[1].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[1].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[1].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[1].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[1].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[1].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[1].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[1].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[1].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[1].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[1].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[1].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[1].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[1].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[1].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[1].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[1].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[1].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[1].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[1].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[1].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[1].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[1].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[1].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[1].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[1].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[1].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[1].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[1].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[1].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[1].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[1].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[1].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[1].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[1].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[1].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[1].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[1].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[1].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[2].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[2].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[2].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[2].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[2].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[2].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[2].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[2].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[2].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[2].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[2].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[2].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[2].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[2].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[2].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[2].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[2].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[2].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[2].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[2].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[2].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[2].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[2].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[2].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[2].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[2].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[2].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[2].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[2].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[2].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[2].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[2].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[2].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[2].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[2].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[2].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[2].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[2].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[2].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[2].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[2].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[2].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[2].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[2].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[2].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[2].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[2].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[2].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[2].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[2].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[2].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[2].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[2].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[2].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[2].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[2].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[2].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[2].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[2].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[2].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[2].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[2].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[2].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[2].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[3].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[3].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[3].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[3].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[3].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[3].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[3].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[3].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[3].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[3].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[3].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[3].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[3].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[3].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[3].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[3].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[3].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[3].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[3].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[3].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[3].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[3].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[3].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[3].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[3].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[3].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[3].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[3].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[3].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[3].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[3].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[3].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[3].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[3].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[3].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[3].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[3].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[3].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[3].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[3].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[3].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[3].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[3].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[3].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[3].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[3].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[3].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[3].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[3].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[3].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[3].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[3].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[3].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[3].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[3].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[3].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[3].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[3].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[3].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[3].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[3].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[3].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[3].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[3].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[4].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[4].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[4].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[4].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[4].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[4].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[4].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[4].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[4].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[4].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[4].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[4].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[4].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[4].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[4].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[4].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[4].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[4].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[4].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[4].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[4].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[4].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[4].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[4].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[4].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[4].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[4].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[4].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[4].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[4].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[4].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[4].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[4].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[4].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[4].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[4].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[4].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[4].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[4].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[4].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[4].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[4].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[4].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[4].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[4].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[4].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[4].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[4].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[4].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[4].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[4].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[4].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[4].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[4].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[4].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[4].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[4].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[4].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[4].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[4].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[4].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[4].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[4].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[4].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[5].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[5].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[5].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[5].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[5].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[5].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[5].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[5].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[5].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[5].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[5].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[5].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[5].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[5].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[5].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[5].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[5].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[5].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[5].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[5].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[5].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[5].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[5].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[5].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[5].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[5].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[5].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[5].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[5].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[5].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[5].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[5].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[5].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[5].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[5].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[5].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[5].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[5].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[5].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[5].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[5].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[5].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[5].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[5].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[5].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[5].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[5].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[5].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[5].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[5].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[5].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[5].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[5].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[5].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[5].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[5].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[5].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[5].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[5].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[5].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[5].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[5].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[5].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[5].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[6].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[6].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[6].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[6].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[6].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[6].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[6].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[6].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[6].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[6].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[6].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[6].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[6].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[6].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[6].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[6].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[6].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[6].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[6].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[6].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[6].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[6].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[6].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[6].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[6].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[6].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[6].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[6].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[6].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[6].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[6].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[6].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[6].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[6].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[6].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[6].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[6].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[6].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[6].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[6].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[6].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[6].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[6].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[6].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[6].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[6].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[6].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[6].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[6].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[6].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[6].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[6].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[6].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[6].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[6].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[6].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[6].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[6].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[6].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[6].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[6].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[6].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[6].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[6].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[7].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[7].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[7].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[7].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[7].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[7].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[7].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[7].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[7].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[7].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[7].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[7].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[7].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[7].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[7].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[7].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[7].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[7].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[7].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[7].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[7].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[7].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[7].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[7].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[7].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[7].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[7].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[7].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[7].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[7].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[7].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[7].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[7].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[7].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[7].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[7].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[7].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[7].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[7].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[7].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[7].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[7].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[7].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[7].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[7].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[7].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[7].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[7].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[7].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[7].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[7].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[7].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[7].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[7].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[7].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[7].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[7].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[7].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[7].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[7].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[7].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[7].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[7].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[7].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[8].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[8].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[8].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[8].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[8].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[8].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[8].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[8].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[8].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[8].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[8].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[8].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[8].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[8].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[8].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[8].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[8].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[8].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[8].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[8].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[8].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[8].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[8].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[8].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[8].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[8].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[8].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[8].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[8].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[8].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[8].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[8].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[8].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[8].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[8].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[8].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[8].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[8].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[8].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[8].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[8].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[8].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[8].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[8].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[8].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[8].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[8].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[8].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[8].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[8].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[8].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[8].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[8].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[8].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[8].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[8].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[8].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[8].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[8].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[8].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[8].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[8].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[8].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[8].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[9].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[9].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[9].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[9].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[9].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[9].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[9].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[9].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[9].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[9].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[9].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[9].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[9].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[9].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[9].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[9].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[9].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[9].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[9].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[9].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[9].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[9].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[9].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[9].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[9].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[9].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[9].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[9].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[9].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[9].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[9].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[9].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[9].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[9].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[9].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[9].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[9].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[9].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[9].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[9].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[9].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[9].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[9].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[9].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[9].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[9].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[9].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[9].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[9].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[9].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[9].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[9].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[9].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[9].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[9].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[9].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[9].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[9].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[9].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[9].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[9].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[9].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[9].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[9].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[10].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[10].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[10].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[10].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[10].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[10].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[10].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[10].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[10].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[10].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[10].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[10].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[10].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[10].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[10].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[10].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[10].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[10].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[10].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[10].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[10].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[10].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[10].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[10].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[10].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[10].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[10].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[10].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[10].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[10].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[10].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[10].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[10].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[10].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[10].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[10].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[10].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[10].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[10].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[10].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[10].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[10].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[10].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[10].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[10].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[10].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[10].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[10].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[10].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[10].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[10].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[10].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[10].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[10].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[10].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[10].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[10].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[10].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[10].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[10].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[10].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[10].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[10].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[10].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[11].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[11].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[11].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[11].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[11].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[11].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[11].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[11].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[11].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[11].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[11].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[11].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[11].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[11].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[11].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[11].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[11].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[11].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[11].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[11].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[11].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[11].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[11].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[11].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[11].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[11].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[11].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[11].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[11].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[11].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[11].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[11].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[11].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[11].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[11].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[11].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[11].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[11].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[11].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[11].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[11].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[11].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[11].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[11].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[11].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[11].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[11].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[11].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[11].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[11].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[11].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[11].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[11].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[11].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[11].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[11].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[11].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[11].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[11].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[11].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[11].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[11].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[11].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[11].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[12].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[12].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[12].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[12].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[12].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[12].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[12].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[12].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[12].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[12].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[12].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[12].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[12].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[12].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[12].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[12].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[12].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[12].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[12].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[12].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[12].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[12].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[12].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[12].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[12].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[12].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[12].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[12].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[12].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[12].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[12].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[12].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[12].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[12].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[12].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[12].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[12].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[12].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[12].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[12].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[12].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[12].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[12].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[12].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[12].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[12].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[12].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[12].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[12].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[12].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[12].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[12].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[12].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[12].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[12].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[12].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[12].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[12].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[12].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[12].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[12].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[12].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[12].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[12].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[13].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[13].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[13].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[13].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[13].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[13].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[13].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[13].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[13].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[13].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[13].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[13].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[13].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[13].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[13].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[13].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[13].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[13].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[13].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[13].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[13].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[13].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[13].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[13].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[13].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[13].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[13].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[13].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[13].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[13].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[13].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[13].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[13].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[13].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[13].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[13].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[13].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[13].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[13].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[13].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[13].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[13].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[13].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[13].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[13].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[13].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[13].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[13].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[13].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[13].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[13].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[13].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[13].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[13].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[13].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[13].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[13].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[13].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[13].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[13].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[13].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[13].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[13].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[13].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[14].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[14].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[14].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[14].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[14].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[14].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[14].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[14].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[14].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[14].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[14].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[14].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[14].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[14].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[14].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[14].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[14].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[14].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[14].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[14].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[14].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[14].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[14].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[14].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[14].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[14].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[14].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[14].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[14].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[14].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[14].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[14].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[14].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[14].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[14].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[14].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[14].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[14].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[14].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[14].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[14].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[14].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[14].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[14].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[14].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[14].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[14].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[14].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[14].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[14].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[14].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[14].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[14].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[14].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[14].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[14].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[14].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[14].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[14].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[14].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[14].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[14].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[14].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[14].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[15].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[15].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[15].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[15].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[15].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[15].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[15].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[15].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[15].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[15].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[15].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[15].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[15].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[15].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[15].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[15].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[15].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[15].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[15].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[15].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[15].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[15].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[15].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[15].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[15].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[15].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[15].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[15].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[15].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[15].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[15].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[15].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[15].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[15].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[15].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[15].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[15].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[15].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[15].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[15].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[15].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[15].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[15].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[15].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[15].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[15].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[15].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[15].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[15].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[15].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[15].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[15].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[15].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[15].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[15].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[15].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[15].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[15].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[15].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[15].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[15].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[15].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[15].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[15].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[16].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[16].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[16].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[16].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[16].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[16].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[16].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[16].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[16].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[16].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[16].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[16].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[16].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[16].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[16].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[16].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[16].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[16].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[16].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[16].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[16].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[16].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[16].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[16].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[16].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[16].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[16].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[16].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[16].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[16].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[16].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[16].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[16].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[16].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[16].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[16].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[16].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[16].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[16].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[16].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[16].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[16].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[16].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[16].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[16].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[16].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[16].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[16].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[16].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[16].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[16].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[16].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[16].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[16].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[16].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[16].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[16].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[16].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[16].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[16].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[16].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[16].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[16].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[16].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[17].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[17].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[17].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[17].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[17].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[17].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[17].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[17].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[17].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[17].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[17].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[17].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[17].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[17].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[17].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[17].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[17].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[17].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[17].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[17].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[17].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[17].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[17].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[17].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[17].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[17].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[17].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[17].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[17].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[17].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[17].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[17].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[17].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[17].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[17].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[17].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[17].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[17].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[17].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[17].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[17].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[17].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[17].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[17].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[17].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[17].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[17].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[17].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[17].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[17].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[17].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[17].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[17].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[17].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[17].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[17].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[17].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[17].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[17].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[17].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[17].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[17].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[17].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[17].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[18].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[18].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[18].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[18].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[18].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[18].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[18].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[18].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[18].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[18].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[18].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[18].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[18].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[18].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[18].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[18].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[18].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[18].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[18].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[18].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[18].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[18].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[18].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[18].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[18].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[18].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[18].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[18].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[18].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[18].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[18].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[18].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[18].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[18].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[18].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[18].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[18].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[18].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[18].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[18].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[18].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[18].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[18].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[18].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[18].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[18].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[18].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[18].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[18].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[18].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[18].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[18].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[18].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[18].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[18].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[18].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[18].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[18].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[18].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[18].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[18].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[18].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[18].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[18].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[19].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[19].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[19].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[19].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[19].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[19].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[19].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[19].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[19].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[19].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[19].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[19].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[19].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[19].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[19].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[19].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[19].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[19].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[19].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[19].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[19].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[19].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[19].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[19].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[19].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[19].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[19].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[19].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[19].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[19].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[19].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[19].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[19].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[19].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[19].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[19].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[19].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[19].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[19].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[19].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[19].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[19].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[19].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[19].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[19].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[19].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[19].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[19].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[19].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[19].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[19].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[19].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[19].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[19].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[19].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[19].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[19].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[19].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[19].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[19].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[19].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[19].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[19].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[19].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[20].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[20].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[20].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[20].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[20].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[20].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[20].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[20].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[20].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[20].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[20].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[20].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[20].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[20].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[20].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[20].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[20].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[20].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[20].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[20].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[20].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[20].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[20].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[20].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[20].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[20].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[20].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[20].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[20].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[20].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[20].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[20].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[20].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[20].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[20].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[20].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[20].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[20].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[20].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[20].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[20].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[20].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[20].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[20].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[20].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[20].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[20].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[20].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[20].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[20].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[20].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[20].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[20].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[20].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[20].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[20].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[20].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[20].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[20].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[20].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[20].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[20].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[20].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[20].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[21].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[21].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[21].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[21].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[21].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[21].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[21].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[21].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[21].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[21].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[21].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[21].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[21].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[21].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[21].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[21].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[21].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[21].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[21].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[21].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[21].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[21].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[21].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[21].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[21].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[21].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[21].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[21].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[21].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[21].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[21].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[21].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[21].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[21].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[21].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[21].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[21].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[21].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[21].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[21].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[21].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[21].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[21].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[21].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[21].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[21].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[21].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[21].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[21].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[21].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[21].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[21].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[21].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[21].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[21].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[21].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[21].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[21].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[21].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[21].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[21].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[21].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[21].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[21].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[22].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[22].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[22].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[22].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[22].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[22].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[22].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[22].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[22].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[22].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[22].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[22].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[22].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[22].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[22].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[22].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[22].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[22].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[22].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[22].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[22].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[22].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[22].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[22].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[22].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[22].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[22].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[22].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[22].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[22].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[22].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[22].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[22].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[22].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[22].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[22].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[22].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[22].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[22].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[22].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[22].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[22].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[22].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[22].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[22].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[22].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[22].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[22].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[22].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[22].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[22].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[22].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[22].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[22].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[22].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[22].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[22].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[22].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[22].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[22].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[22].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[22].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[22].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[22].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[23].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[23].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[23].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[23].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[23].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[23].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[23].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[23].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[23].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[23].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[23].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[23].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[23].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[23].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[23].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[23].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[23].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[23].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[23].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[23].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[23].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[23].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[23].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[23].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[23].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[23].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[23].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[23].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[23].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[23].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[23].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[23].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[23].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[23].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[23].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[23].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[23].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[23].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[23].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[23].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[23].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[23].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[23].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[23].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[23].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[23].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[23].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[23].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[23].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[23].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[23].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[23].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[23].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[23].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[23].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[23].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[23].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[23].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[23].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[23].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[23].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[23].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[23].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[23].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[24].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[24].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[24].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[24].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[24].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[24].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[24].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[24].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[24].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[24].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[24].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[24].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[24].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[24].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[24].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[24].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[24].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[24].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[24].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[24].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[24].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[24].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[24].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[24].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[24].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[24].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[24].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[24].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[24].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[24].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[24].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[24].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[24].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[24].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[24].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[24].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[24].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[24].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[24].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[24].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[24].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[24].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[24].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[24].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[24].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[24].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[24].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[24].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[24].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[24].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[24].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[24].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[24].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[24].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[24].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[24].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[24].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[24].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[24].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[24].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[24].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[24].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[24].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[24].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[25].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[25].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[25].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[25].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[25].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[25].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[25].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[25].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[25].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[25].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[25].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[25].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[25].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[25].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[25].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[25].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[25].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[25].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[25].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[25].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[25].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[25].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[25].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[25].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[25].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[25].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[25].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[25].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[25].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[25].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[25].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[25].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[25].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[25].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[25].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[25].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[25].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[25].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[25].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[25].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[25].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[25].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[25].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[25].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[25].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[25].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[25].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[25].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[25].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[25].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[25].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[25].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[25].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[25].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[25].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[25].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[25].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[25].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[25].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[25].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[25].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[25].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[25].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[25].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[26].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[26].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[26].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[26].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[26].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[26].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[26].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[26].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[26].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[26].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[26].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[26].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[26].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[26].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[26].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[26].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[26].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[26].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[26].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[26].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[26].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[26].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[26].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[26].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[26].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[26].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[26].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[26].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[26].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[26].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[26].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[26].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[26].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[26].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[26].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[26].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[26].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[26].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[26].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[26].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[26].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[26].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[26].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[26].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[26].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[26].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[26].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[26].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[26].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[26].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[26].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[26].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[26].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[26].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[26].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[26].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[26].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[26].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[26].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[26].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[26].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[26].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[26].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[26].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[27].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[27].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[27].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[27].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[27].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[27].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[27].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[27].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[27].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[27].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[27].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[27].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[27].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[27].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[27].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[27].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[27].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[27].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[27].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[27].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[27].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[27].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[27].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[27].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[27].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[27].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[27].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[27].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[27].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[27].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[27].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[27].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[27].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[27].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[27].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[27].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[27].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[27].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[27].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[27].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[27].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[27].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[27].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[27].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[27].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[27].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[27].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[27].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[27].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[27].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[27].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[27].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[27].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[27].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[27].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[27].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[27].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[27].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[27].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[27].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[27].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[27].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[27].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[27].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[28].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[28].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[28].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[28].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[28].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[28].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[28].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[28].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[28].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[28].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[28].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[28].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[28].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[28].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[28].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[28].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[28].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[28].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[28].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[28].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[28].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[28].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[28].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[28].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[28].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[28].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[28].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[28].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[28].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[28].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[28].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[28].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[28].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[28].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[28].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[28].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[28].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[28].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[28].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[28].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[28].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[28].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[28].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[28].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[28].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[28].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[28].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[28].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[28].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[28].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[28].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[28].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[28].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[28].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[28].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[28].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[28].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[28].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[28].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[28].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[28].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[28].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[28].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[28].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[29].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[29].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[29].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[29].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[29].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[29].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[29].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[29].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[29].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[29].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[29].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[29].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[29].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[29].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[29].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[29].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[29].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[29].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[29].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[29].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[29].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[29].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[29].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[29].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[29].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[29].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[29].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[29].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[29].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[29].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[29].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[29].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[29].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[29].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[29].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[29].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[29].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[29].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[29].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[29].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[29].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[29].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[29].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[29].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[29].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[29].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[29].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[29].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[29].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[29].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[29].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[29].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[29].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[29].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[29].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[29].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[29].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[29].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[29].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[29].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[29].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[29].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[29].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[29].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[30].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[30].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[30].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[30].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[30].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[30].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[30].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[30].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[30].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[30].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[30].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[30].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[30].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[30].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[30].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[30].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[30].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[30].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[30].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[30].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[30].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[30].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[30].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[30].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[30].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[30].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[30].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[30].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[30].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[30].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[30].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[30].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[30].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[30].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[30].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[30].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[30].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[30].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[30].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[30].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[30].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[30].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[30].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[30].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[30].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[30].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[30].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[30].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[30].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[30].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[30].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[30].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[30].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[30].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[30].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[30].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[30].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[30].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[30].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[30].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[30].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[30].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[30].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[30].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[31].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[31].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[31].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[31].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[31].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[31].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[31].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[31].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[31].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[31].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[31].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[31].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[31].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[31].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[31].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[31].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[31].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[31].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[31].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[31].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[31].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[31].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[31].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[31].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[31].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[31].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[31].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[31].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[31].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[31].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[31].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[31].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[31].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[31].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[31].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[31].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[31].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[31].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[31].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[31].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[31].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[31].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[31].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[31].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[31].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[31].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[31].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[31].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[31].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[31].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[31].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[31].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[31].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[31].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[31].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[31].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[31].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[31].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[31].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[31].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[31].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[31].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[31].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[31].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[32].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[32].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[32].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[32].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[32].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[32].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[32].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[32].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[32].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[32].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[32].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[32].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[32].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[32].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[32].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[32].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[32].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[32].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[32].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[32].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[32].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[32].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[32].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[32].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[32].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[32].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[32].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[32].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[32].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[32].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[32].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[32].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[32].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[32].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[32].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[32].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[32].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[32].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[32].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[32].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[32].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[32].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[32].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[32].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[32].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[32].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[32].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[32].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[32].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[32].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[32].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[32].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[32].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[32].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[32].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[32].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[32].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[32].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[32].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[32].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[32].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[32].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[32].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[32].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[33].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[33].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[33].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[33].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[33].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[33].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[33].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[33].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[33].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[33].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[33].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[33].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[33].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[33].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[33].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[33].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[33].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[33].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[33].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[33].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[33].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[33].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[33].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[33].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[33].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[33].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[33].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[33].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[33].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[33].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[33].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[33].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[33].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[33].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[33].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[33].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[33].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[33].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[33].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[33].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[33].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[33].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[33].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[33].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[33].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[33].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[33].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[33].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[33].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[33].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[33].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[33].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[33].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[33].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[33].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[33].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[33].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[33].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[33].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[33].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[33].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[33].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[33].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[33].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[34].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[34].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[34].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[34].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[34].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[34].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[34].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[34].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[34].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[34].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[34].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[34].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[34].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[34].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[34].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[34].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[34].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[34].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[34].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[34].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[34].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[34].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[34].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[34].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[34].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[34].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[34].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[34].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[34].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[34].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[34].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[34].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[34].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[34].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[34].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[34].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[34].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[34].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[34].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[34].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[34].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[34].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[34].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[34].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[34].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[34].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[34].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[34].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[34].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[34].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[34].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[34].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[34].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[34].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[34].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[34].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[34].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[34].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[34].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[34].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[34].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[34].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[34].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[34].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[35].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[35].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[35].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[35].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[35].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[35].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[35].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[35].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[35].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[35].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[35].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[35].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[35].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[35].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[35].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[35].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[35].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[35].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[35].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[35].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[35].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[35].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[35].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[35].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[35].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[35].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[35].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[35].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[35].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[35].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[35].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[35].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[35].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[35].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[35].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[35].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[35].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[35].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[35].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[35].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[35].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[35].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[35].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[35].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[35].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[35].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[35].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[35].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[35].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[35].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[35].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[35].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[35].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[35].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[35].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[35].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[35].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[35].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[35].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[35].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[35].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[35].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[35].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[35].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[36].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[36].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[36].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[36].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[36].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[36].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[36].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[36].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[36].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[36].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[36].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[36].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[36].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[36].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[36].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[36].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[36].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[36].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[36].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[36].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[36].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[36].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[36].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[36].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[36].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[36].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[36].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[36].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[36].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[36].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[36].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[36].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[36].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[36].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[36].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[36].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[36].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[36].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[36].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[36].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[36].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[36].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[36].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[36].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[36].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[36].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[36].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[36].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[36].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[36].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[36].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[36].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[36].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[36].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[36].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[36].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[36].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[36].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[36].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[36].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[36].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[36].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[36].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[36].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[37].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[37].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[37].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[37].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[37].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[37].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[37].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[37].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[37].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[37].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[37].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[37].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[37].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[37].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[37].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[37].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[37].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[37].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[37].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[37].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[37].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[37].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[37].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[37].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[37].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[37].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[37].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[37].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[37].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[37].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[37].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[37].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[37].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[37].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[37].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[37].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[37].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[37].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[37].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[37].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[37].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[37].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[37].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[37].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[37].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[37].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[37].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[37].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[37].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[37].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[37].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[37].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[37].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[37].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[37].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[37].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[37].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[37].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[37].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[37].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[37].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[37].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[37].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[37].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[38].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[38].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[38].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[38].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[38].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[38].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[38].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[38].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[38].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[38].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[38].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[38].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[38].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[38].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[38].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[38].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[38].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[38].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[38].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[38].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[38].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[38].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[38].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[38].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[38].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[38].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[38].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[38].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[38].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[38].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[38].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[38].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[38].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[38].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[38].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[38].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[38].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[38].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[38].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[38].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[38].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[38].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[38].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[38].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[38].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[38].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[38].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[38].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[38].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[38].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[38].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[38].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[38].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[38].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[38].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[38].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[38].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[38].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[38].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[38].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[38].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[38].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[38].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[38].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[39].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[39].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[39].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[39].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[39].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[39].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[39].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[39].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[39].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[39].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[39].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[39].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[39].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[39].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[39].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[39].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[39].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[39].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[39].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[39].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[39].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[39].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[39].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[39].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[39].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[39].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[39].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[39].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[39].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[39].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[39].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[39].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[39].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[39].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[39].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[39].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[39].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[39].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[39].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[39].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[39].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[39].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[39].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[39].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[39].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[39].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[39].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[39].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[39].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[39].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[39].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[39].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[39].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[39].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[39].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[39].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[39].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[39].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[39].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[39].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[39].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[39].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[39].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[39].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[40].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[40].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[40].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[40].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[40].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[40].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[40].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[40].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[40].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[40].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[40].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[40].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[40].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[40].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[40].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[40].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[40].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[40].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[40].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[40].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[40].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[40].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[40].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[40].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[40].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[40].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[40].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[40].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[40].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[40].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[40].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[40].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[40].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[40].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[40].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[40].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[40].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[40].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[40].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[40].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[40].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[40].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[40].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[40].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[40].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[40].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[40].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[40].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[40].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[40].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[40].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[40].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[40].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[40].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[40].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[40].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[40].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[40].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[40].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[40].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[40].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[40].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[40].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[40].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[41].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[41].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[41].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[41].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[41].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[41].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[41].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[41].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[41].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[41].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[41].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[41].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[41].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[41].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[41].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[41].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[41].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[41].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[41].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[41].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[41].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[41].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[41].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[41].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[41].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[41].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[41].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[41].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[41].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[41].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[41].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[41].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[41].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[41].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[41].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[41].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[41].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[41].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[41].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[41].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[41].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[41].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[41].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[41].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[41].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[41].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[41].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[41].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[41].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[41].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[41].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[41].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[41].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[41].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[41].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[41].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[41].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[41].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[41].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[41].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[41].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[41].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[41].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[41].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[42].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[42].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[42].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[42].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[42].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[42].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[42].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[42].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[42].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[42].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[42].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[42].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[42].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[42].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[42].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[42].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[42].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[42].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[42].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[42].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[42].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[42].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[42].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[42].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[42].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[42].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[42].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[42].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[42].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[42].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[42].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[42].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[42].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[42].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[42].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[42].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[42].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[42].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[42].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[42].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[42].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[42].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[42].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[42].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[42].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[42].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[42].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[42].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[42].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[42].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[42].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[42].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[42].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[42].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[42].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[42].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[42].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[42].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[42].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[42].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[42].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[42].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[42].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[42].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[43].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[43].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[43].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[43].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[43].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[43].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[43].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[43].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[43].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[43].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[43].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[43].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[43].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[43].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[43].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[43].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[43].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[43].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[43].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[43].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[43].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[43].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[43].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[43].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[43].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[43].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[43].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[43].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[43].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[43].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[43].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[43].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[43].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[43].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[43].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[43].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[43].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[43].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[43].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[43].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[43].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[43].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[43].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[43].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[43].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[43].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[43].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[43].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[43].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[43].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[43].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[43].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[43].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[43].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[43].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[43].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[43].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[43].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[43].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[43].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[43].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[43].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[43].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[43].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[44].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[44].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[44].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[44].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[44].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[44].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[44].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[44].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[44].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[44].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[44].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[44].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[44].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[44].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[44].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[44].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[44].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[44].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[44].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[44].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[44].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[44].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[44].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[44].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[44].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[44].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[44].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[44].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[44].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[44].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[44].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[44].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[44].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[44].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[44].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[44].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[44].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[44].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[44].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[44].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[44].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[44].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[44].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[44].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[44].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[44].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[44].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[44].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[44].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[44].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[44].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[44].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[44].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[44].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[44].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[44].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[44].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[44].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[44].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[44].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[44].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[44].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[44].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[44].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[45].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[45].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[45].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[45].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[45].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[45].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[45].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[45].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[45].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[45].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[45].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[45].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[45].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[45].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[45].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[45].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[45].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[45].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[45].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[45].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[45].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[45].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[45].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[45].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[45].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[45].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[45].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[45].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[45].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[45].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[45].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[45].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[45].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[45].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[45].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[45].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[45].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[45].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[45].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[45].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[45].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[45].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[45].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[45].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[45].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[45].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[45].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[45].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[45].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[45].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[45].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[45].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[45].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[45].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[45].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[45].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[45].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[45].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[45].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[45].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[45].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[45].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[45].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[45].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[46].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[46].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[46].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[46].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[46].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[46].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[46].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[46].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[46].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[46].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[46].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[46].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[46].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[46].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[46].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[46].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[46].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[46].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[46].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[46].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[46].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[46].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[46].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[46].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[46].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[46].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[46].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[46].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[46].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[46].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[46].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[46].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[46].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[46].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[46].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[46].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[46].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[46].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[46].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[46].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[46].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[46].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[46].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[46].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[46].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[46].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[46].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[46].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[46].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[46].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[46].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[46].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[46].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[46].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[46].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[46].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[46].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[46].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[46].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[46].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[46].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[46].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[46].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[46].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[47].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[47].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[47].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[47].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[47].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[47].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[47].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[47].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[47].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[47].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[47].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[47].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[47].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[47].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[47].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[47].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[47].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[47].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[47].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[47].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[47].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[47].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[47].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[47].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[47].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[47].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[47].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[47].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[47].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[47].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[47].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[47].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[47].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[47].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[47].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[47].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[47].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[47].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[47].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[47].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[47].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[47].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[47].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[47].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[47].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[47].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[47].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[47].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[47].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[47].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[47].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[47].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[47].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[47].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[47].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[47].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[47].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[47].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[47].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[47].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[47].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[47].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[47].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[47].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[48].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[48].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[48].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[48].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[48].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[48].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[48].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[48].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[48].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[48].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[48].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[48].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[48].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[48].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[48].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[48].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[48].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[48].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[48].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[48].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[48].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[48].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[48].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[48].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[48].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[48].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[48].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[48].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[48].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[48].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[48].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[48].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[48].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[48].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[48].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[48].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[48].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[48].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[48].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[48].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[48].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[48].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[48].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[48].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[48].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[48].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[48].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[48].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[48].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[48].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[48].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[48].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[48].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[48].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[48].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[48].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[48].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[48].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[48].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[48].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[48].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[48].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[48].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[48].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[49].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[49].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[49].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[49].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[49].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[49].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[49].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[49].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[49].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[49].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[49].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[49].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[49].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[49].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[49].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[49].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[49].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[49].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[49].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[49].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[49].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[49].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[49].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[49].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[49].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[49].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[49].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[49].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[49].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[49].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[49].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[49].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[49].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[49].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[49].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[49].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[49].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[49].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[49].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[49].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[49].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[49].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[49].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[49].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[49].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[49].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[49].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[49].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[49].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[49].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[49].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[49].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[49].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[49].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[49].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[49].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[49].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[49].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[49].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[49].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[49].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[49].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[49].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[49].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[50].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[50].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[50].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[50].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[50].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[50].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[50].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[50].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[50].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[50].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[50].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[50].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[50].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[50].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[50].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[50].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[50].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[50].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[50].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[50].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[50].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[50].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[50].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[50].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[50].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[50].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[50].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[50].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[50].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[50].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[50].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[50].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[50].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[50].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[50].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[50].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[50].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[50].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[50].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[50].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[50].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[50].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[50].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[50].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[50].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[50].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[50].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[50].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[50].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[50].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[50].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[50].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[50].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[50].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[50].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[50].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[50].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[50].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[50].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[50].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[50].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[50].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[50].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[50].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[51].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[51].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[51].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[51].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[51].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[51].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[51].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[51].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[51].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[51].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[51].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[51].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[51].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[51].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[51].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[51].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[51].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[51].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[51].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[51].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[51].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[51].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[51].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[51].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[51].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[51].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[51].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[51].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[51].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[51].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[51].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[51].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[51].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[51].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[51].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[51].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[51].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[51].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[51].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[51].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[51].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[51].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[51].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[51].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[51].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[51].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[51].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[51].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[51].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[51].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[51].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[51].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[51].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[51].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[51].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[51].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[51].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[51].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[51].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[51].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[51].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[51].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[51].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[51].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[52].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[52].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[52].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[52].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[52].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[52].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[52].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[52].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[52].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[52].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[52].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[52].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[52].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[52].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[52].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[52].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[52].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[52].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[52].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[52].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[52].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[52].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[52].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[52].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[52].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[52].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[52].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[52].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[52].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[52].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[52].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[52].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[52].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[52].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[52].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[52].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[52].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[52].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[52].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[52].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[52].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[52].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[52].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[52].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[52].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[52].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[52].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[52].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[52].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[52].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[52].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[52].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[52].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[52].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[52].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[52].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[52].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[52].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[52].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[52].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[52].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[52].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[52].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[52].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[53].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[53].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[53].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[53].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[53].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[53].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[53].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[53].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[53].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[53].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[53].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[53].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[53].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[53].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[53].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[53].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[53].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[53].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[53].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[53].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[53].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[53].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[53].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[53].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[53].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[53].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[53].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[53].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[53].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[53].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[53].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[53].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[53].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[53].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[53].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[53].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[53].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[53].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[53].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[53].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[53].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[53].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[53].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[53].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[53].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[53].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[53].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[53].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[53].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[53].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[53].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[53].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[53].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[53].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[53].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[53].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[53].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[53].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[53].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[53].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[53].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[53].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[53].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[53].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[54].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[54].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[54].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[54].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[54].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[54].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[54].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[54].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[54].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[54].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[54].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[54].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[54].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[54].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[54].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[54].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[54].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[54].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[54].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[54].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[54].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[54].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[54].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[54].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[54].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[54].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[54].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[54].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[54].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[54].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[54].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[54].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[54].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[54].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[54].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[54].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[54].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[54].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[54].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[54].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[54].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[54].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[54].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[54].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[54].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[54].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[54].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[54].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[54].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[54].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[54].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[54].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[54].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[54].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[54].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[54].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[54].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[54].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[54].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[54].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[54].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[54].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[54].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[54].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[55].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[55].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[55].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[55].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[55].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[55].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[55].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[55].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[55].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[55].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[55].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[55].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[55].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[55].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[55].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[55].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[55].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[55].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[55].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[55].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[55].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[55].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[55].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[55].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[55].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[55].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[55].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[55].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[55].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[55].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[55].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[55].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[55].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[55].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[55].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[55].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[55].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[55].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[55].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[55].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[55].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[55].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[55].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[55].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[55].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[55].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[55].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[55].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[55].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[55].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[55].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[55].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[55].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[55].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[55].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[55].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[55].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[55].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[55].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[55].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[55].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[55].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[55].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[55].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[56].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[56].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[56].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[56].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[56].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[56].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[56].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[56].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[56].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[56].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[56].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[56].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[56].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[56].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[56].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[56].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[56].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[56].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[56].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[56].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[56].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[56].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[56].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[56].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[56].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[56].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[56].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[56].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[56].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[56].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[56].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[56].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[56].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[56].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[56].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[56].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[56].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[56].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[56].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[56].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[56].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[56].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[56].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[56].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[56].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[56].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[56].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[56].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[56].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[56].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[56].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[56].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[56].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[56].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[56].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[56].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[56].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[56].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[56].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[56].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[56].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[56].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[56].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[56].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[57].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[57].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[57].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[57].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[57].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[57].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[57].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[57].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[57].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[57].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[57].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[57].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[57].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[57].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[57].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[57].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[57].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[57].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[57].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[57].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[57].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[57].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[57].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[57].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[57].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[57].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[57].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[57].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[57].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[57].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[57].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[57].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[57].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[57].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[57].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[57].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[57].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[57].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[57].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[57].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[57].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[57].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[57].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[57].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[57].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[57].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[57].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[57].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[57].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[57].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[57].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[57].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[57].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[57].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[57].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[57].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[57].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[57].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[57].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[57].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[57].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[57].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[57].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[57].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[58].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[58].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[58].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[58].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[58].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[58].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[58].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[58].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[58].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[58].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[58].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[58].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[58].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[58].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[58].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[58].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[58].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[58].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[58].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[58].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[58].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[58].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[58].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[58].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[58].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[58].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[58].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[58].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[58].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[58].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[58].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[58].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[58].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[58].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[58].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[58].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[58].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[58].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[58].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[58].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[58].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[58].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[58].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[58].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[58].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[58].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[58].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[58].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[58].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[58].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[58].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[58].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[58].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[58].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[58].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[58].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[58].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[58].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[58].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[58].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[58].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[58].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[58].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[58].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[59].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[59].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[59].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[59].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[59].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[59].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[59].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[59].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[59].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[59].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[59].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[59].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[59].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[59].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[59].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[59].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[59].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[59].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[59].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[59].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[59].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[59].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[59].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[59].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[59].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[59].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[59].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[59].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[59].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[59].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[59].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[59].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[59].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[59].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[59].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[59].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[59].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[59].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[59].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[59].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[59].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[59].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[59].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[59].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[59].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[59].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[59].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[59].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[59].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[59].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[59].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[59].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[59].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[59].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[59].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[59].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[59].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[59].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[59].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[59].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[59].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[59].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[59].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[59].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[60].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[60].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[60].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[60].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[60].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[60].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[60].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[60].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[60].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[60].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[60].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[60].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[60].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[60].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[60].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[60].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[60].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[60].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[60].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[60].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[60].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[60].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[60].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[60].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[60].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[60].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[60].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[60].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[60].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[60].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[60].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[60].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[60].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[60].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[60].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[60].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[60].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[60].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[60].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[60].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[60].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[60].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[60].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[60].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[60].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[60].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[60].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[60].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[60].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[60].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[60].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[60].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[60].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[60].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[60].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[60].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[60].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[60].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[60].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[60].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[60].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[60].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[60].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[60].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[61].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[61].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[61].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[61].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[61].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[61].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[61].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[61].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[61].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[61].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[61].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[61].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[61].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[61].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[61].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[61].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[61].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[61].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[61].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[61].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[61].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[61].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[61].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[61].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[61].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[61].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[61].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[61].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[61].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[61].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[61].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[61].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[61].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[61].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[61].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[61].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[61].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[61].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[61].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[61].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[61].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[61].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[61].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[61].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[61].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[61].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[61].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[61].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[61].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[61].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[61].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[61].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[61].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[61].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[61].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[61].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[61].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[61].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[61].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[61].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[61].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[61].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[61].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[61].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[62].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[62].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[62].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[62].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[62].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[62].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[62].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[62].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[62].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[62].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[62].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[62].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[62].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[62].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[62].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[62].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[62].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[62].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[62].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[62].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[62].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[62].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[62].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[62].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[62].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[62].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[62].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[62].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[62].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[62].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[62].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[62].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[62].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[62].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[62].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[62].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[62].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[62].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[62].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[62].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[62].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[62].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[62].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[62].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[62].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[62].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[62].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[62].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[62].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[62].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[62].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[62].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[62].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[62].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[62].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[62].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[62].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[62].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[62].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[62].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[62].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[62].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[62].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[62].pe.lane31_r135 = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[63].pe.lane0_r134 = 32'h0010;
            force pe_array_inst.pe_inst[63].pe.lane1_r134 = 32'h1010;
            force pe_array_inst.pe_inst[63].pe.lane2_r134 = 32'h2010;
            force pe_array_inst.pe_inst[63].pe.lane3_r134 = 32'h3010;
            force pe_array_inst.pe_inst[63].pe.lane4_r134 = 32'h4010;
            force pe_array_inst.pe_inst[63].pe.lane5_r134 = 32'h5010;
            force pe_array_inst.pe_inst[63].pe.lane6_r134 = 32'h6010;
            force pe_array_inst.pe_inst[63].pe.lane7_r134 = 32'h7010;
            force pe_array_inst.pe_inst[63].pe.lane8_r134 = 32'h8010;
            force pe_array_inst.pe_inst[63].pe.lane9_r134 = 32'h9010;
            force pe_array_inst.pe_inst[63].pe.lane10_r134 = 32'ha010;
            force pe_array_inst.pe_inst[63].pe.lane11_r134 = 32'hb010;
            force pe_array_inst.pe_inst[63].pe.lane12_r134 = 32'hc010;
            force pe_array_inst.pe_inst[63].pe.lane13_r134 = 32'hd010;
            force pe_array_inst.pe_inst[63].pe.lane14_r134 = 32'he010;
            force pe_array_inst.pe_inst[63].pe.lane15_r134 = 32'hf010;
            force pe_array_inst.pe_inst[63].pe.lane16_r134 = 32'h10010;
            force pe_array_inst.pe_inst[63].pe.lane17_r134 = 32'h11010;
            force pe_array_inst.pe_inst[63].pe.lane18_r134 = 32'h12010;
            force pe_array_inst.pe_inst[63].pe.lane19_r134 = 32'h13010;
            force pe_array_inst.pe_inst[63].pe.lane20_r134 = 32'h14010;
            force pe_array_inst.pe_inst[63].pe.lane21_r134 = 32'h15010;
            force pe_array_inst.pe_inst[63].pe.lane22_r134 = 32'h16010;
            force pe_array_inst.pe_inst[63].pe.lane23_r134 = 32'h17010;
            force pe_array_inst.pe_inst[63].pe.lane24_r134 = 32'h18010;
            force pe_array_inst.pe_inst[63].pe.lane25_r134 = 32'h19010;
            force pe_array_inst.pe_inst[63].pe.lane26_r134 = 32'h1a010;
            force pe_array_inst.pe_inst[63].pe.lane27_r134 = 32'h1b010;
            force pe_array_inst.pe_inst[63].pe.lane28_r134 = 32'h1c010;
            force pe_array_inst.pe_inst[63].pe.lane29_r134 = 32'h1d010;
            force pe_array_inst.pe_inst[63].pe.lane30_r134 = 32'h1e010;
            force pe_array_inst.pe_inst[63].pe.lane31_r134 = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[63].pe.lane0_r135 = 32'h0800;
            force pe_array_inst.pe_inst[63].pe.lane1_r135 = 32'h1800;
            force pe_array_inst.pe_inst[63].pe.lane2_r135 = 32'h2800;
            force pe_array_inst.pe_inst[63].pe.lane3_r135 = 32'h3800;
            force pe_array_inst.pe_inst[63].pe.lane4_r135 = 32'h4800;
            force pe_array_inst.pe_inst[63].pe.lane5_r135 = 32'h5800;
            force pe_array_inst.pe_inst[63].pe.lane6_r135 = 32'h6800;
            force pe_array_inst.pe_inst[63].pe.lane7_r135 = 32'h7800;
            force pe_array_inst.pe_inst[63].pe.lane8_r135 = 32'h8800;
            force pe_array_inst.pe_inst[63].pe.lane9_r135 = 32'h9800;
            force pe_array_inst.pe_inst[63].pe.lane10_r135 = 32'ha800;
            force pe_array_inst.pe_inst[63].pe.lane11_r135 = 32'hb800;
            force pe_array_inst.pe_inst[63].pe.lane12_r135 = 32'hc800;
            force pe_array_inst.pe_inst[63].pe.lane13_r135 = 32'hd800;
            force pe_array_inst.pe_inst[63].pe.lane14_r135 = 32'he800;
            force pe_array_inst.pe_inst[63].pe.lane15_r135 = 32'hf800;
            force pe_array_inst.pe_inst[63].pe.lane16_r135 = 32'h10800;
            force pe_array_inst.pe_inst[63].pe.lane17_r135 = 32'h11800;
            force pe_array_inst.pe_inst[63].pe.lane18_r135 = 32'h12800;
            force pe_array_inst.pe_inst[63].pe.lane19_r135 = 32'h13800;
            force pe_array_inst.pe_inst[63].pe.lane20_r135 = 32'h14800;
            force pe_array_inst.pe_inst[63].pe.lane21_r135 = 32'h15800;
            force pe_array_inst.pe_inst[63].pe.lane22_r135 = 32'h16800;
            force pe_array_inst.pe_inst[63].pe.lane23_r135 = 32'h17800;
            force pe_array_inst.pe_inst[63].pe.lane24_r135 = 32'h18800;
            force pe_array_inst.pe_inst[63].pe.lane25_r135 = 32'h19800;
            force pe_array_inst.pe_inst[63].pe.lane26_r135 = 32'h1a800;
            force pe_array_inst.pe_inst[63].pe.lane27_r135 = 32'h1b800;
            force pe_array_inst.pe_inst[63].pe.lane28_r135 = 32'h1c800;
            force pe_array_inst.pe_inst[63].pe.lane29_r135 = 32'h1d800;
            force pe_array_inst.pe_inst[63].pe.lane30_r135 = 32'h1e800;
            force pe_array_inst.pe_inst[63].pe.lane31_r135 = 32'h1f800;

            // ##################################################
            // DMA Type and length of stream

            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[0].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[0].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[1].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[1].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[2].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[2].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[3].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[3].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[4].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[4].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[4].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[4].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[5].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[5].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[5].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[5].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[6].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[6].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[6].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[6].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[7].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[7].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[7].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[7].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[8].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[8].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[8].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[8].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[9].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[9].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[9].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[9].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[10].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[10].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[10].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[10].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[11].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[11].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[11].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[11].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[12].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[12].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[12].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[12].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[13].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[13].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[13].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[13].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[14].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[14].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[14].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[14].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[15].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[15].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[15].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[15].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[16].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[16].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[16].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[16].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[17].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[17].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[17].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[17].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[18].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[18].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[18].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[18].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[19].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[19].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[19].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[19].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[20].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[20].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[20].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[20].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[21].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[21].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[21].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[21].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[22].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[22].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[22].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[22].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[23].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[23].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[23].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[23].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[24].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[24].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[24].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[24].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[25].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[25].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[25].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[25].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[26].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[26].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[26].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[26].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[27].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[27].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[27].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[27].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[28].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[28].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[28].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[28].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[29].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[29].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[29].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[29].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[30].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[30].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[30].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[30].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[31].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[31].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[31].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[31].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[32].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[32].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[32].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[32].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[33].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[33].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[33].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[33].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[34].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[34].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[34].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[34].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[35].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[35].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[35].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[35].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[36].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[36].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[36].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[36].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[37].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[37].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[37].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[37].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[38].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[38].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[38].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[38].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[39].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[39].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[39].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[39].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[40].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[40].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[40].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[40].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[41].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[41].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[41].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[41].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[42].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[42].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[42].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[42].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[43].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[43].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[43].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[43].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[44].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[44].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[44].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[44].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[45].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[45].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[45].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[45].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[46].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[46].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[46].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[46].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[47].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[47].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[47].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[47].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[48].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[48].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[48].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[48].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[49].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[49].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[49].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[49].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[50].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[50].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[50].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[50].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[51].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[51].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[51].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[51].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[52].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[52].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[52].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[52].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[53].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[53].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[53].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[53].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[54].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[54].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[54].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[54].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[55].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[55].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[55].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[55].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[56].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[56].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[56].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[56].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[57].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[57].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[57].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[57].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[58].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[58].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[58].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[58].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[59].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[59].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[59].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[59].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[60].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[60].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[60].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[60].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[61].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[61].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[61].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[61].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[62].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[62].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[62].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[62].pe.lane31_r133[15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[63].pe.lane0_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane0_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane1_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane1_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane2_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane2_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane3_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane3_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane4_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane4_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane5_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane5_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane6_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane6_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane7_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane7_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane8_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane8_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane9_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane9_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane10_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane10_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane11_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane11_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane12_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane12_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane13_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane13_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane14_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane14_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane15_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane15_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane16_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane16_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane17_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane17_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane18_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane18_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane19_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane19_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane20_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane20_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane21_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane21_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane22_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane22_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane23_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane23_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane24_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane24_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane25_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane25_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane26_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane26_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane27_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane27_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane28_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane28_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane29_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane29_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane30_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane30_r132[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane31_r132[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane31_r132[15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[63].pe.lane0_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane0_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane1_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane1_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane2_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane2_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane3_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane3_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane4_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane4_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane5_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane5_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane6_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane6_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane7_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane7_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane8_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane8_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane9_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane9_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane10_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane10_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane11_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane11_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane12_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane12_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane13_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane13_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane14_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane14_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane15_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane15_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane16_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane16_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane17_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane17_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane18_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane18_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane19_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane19_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane20_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane20_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane21_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane21_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane22_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane22_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane23_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane23_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane24_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane24_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane25_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane25_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane26_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane26_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane27_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane27_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane28_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane28_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane29_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane29_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane30_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane30_r133[15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[63].pe.lane31_r133[19:16] = 4'd4;
            force pe_array_inst.pe_inst[63].pe.lane31_r133[15:0]  = numOfTypes;

            // ##################################################
            // Enable and set transfer type

            repeat(10) @(negedge clk); 

            // Enable
            force pe_array_inst.pe_inst[0].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[1].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[2].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[3].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[4].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[5].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[6].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[7].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[8].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[9].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[10].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[11].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[12].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[13].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[14].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[15].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[16].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[17].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[18].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[19].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[20].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[21].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[22].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[23].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[24].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[25].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[26].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[27].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[28].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[29].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[30].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[31].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[32].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[33].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[34].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[35].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[36].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[37].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[38].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[39].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[40].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[41].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[42].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[43].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[44].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[45].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[46].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[47].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[48].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[49].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[50].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[51].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[52].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[53].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[54].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[55].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[56].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[57].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[58].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[59].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[60].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[61].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[62].pe.rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[63].pe.rs0[0]           = 1'b1;

            // Operation
            force pe_array_inst.pe_inst[0].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[1].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[2].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[3].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[4].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[5].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[6].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[7].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[8].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[9].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[10].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[11].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[12].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[13].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[14].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[15].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[16].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[17].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[18].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[19].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[20].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[21].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[22].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[23].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[24].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[25].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[26].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[27].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[28].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[29].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[30].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[31].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[32].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[33].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[34].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[35].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[36].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[37].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[38].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[39].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[40].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[41].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[42].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[43].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[44].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[45].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[46].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[47].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[48].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[49].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[50].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[51].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[52].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[53].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[54].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[55].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[56].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[57].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[58].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[59].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[60].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[61].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[62].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[63].pe.rs0[15:1] = `STREAMING_OP_CNTL_OPERATION_FP_MAC_FROM_EXT_TO_MEM ;

            repeat(50) @(negedge clk);