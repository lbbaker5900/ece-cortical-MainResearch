/*****************************************************************

    File name   : noc_cntl.vh
    Author      : Lee Baker
    Affiliation : North Carolina State University, Raleigh, NC
    Date        : Aug 2015
    email       : lbbaker@ncsu.edu

*****************************************************************/

`define NOC_CONT_EXTERNAL_DATA_WIDTH         42
`define NOC_CONT_EXTERNAL_DATA_MSB           `NOC_CONT_EXTERNAL_DATA_WIDTH-1
`define NOC_CONT_EXTERNAL_DATA_LSB           0
`define NOC_CONT_EXTERNAL_DATA_RANGE         `NOC_CONT_EXTERNAL_DATA_MSB : `NOC_CONT_EXTERNAL_DATA_LSB

`define NOC_CONT_INTERNAL_DATA_WIDTH         `PE_NOC_INTERNAL_DATA_WIDTH
`define NOC_CONT_INTERNAL_DATA_MSB           `NOC_CONT_INTERNAL_DATA_WIDTH-1
`define NOC_CONT_INTERNAL_DATA_LSB           0
`define NOC_CONT_INTERNAL_DATA_RANGE         `NOC_CONT_INTERNAL_DATA_MSB : `NOC_CONT_INTERNAL_DATA_LSB

`define NOC_CONT_EXT_DATA_TO_INT_DATA_RANGE         `PE_EXEC_LANE_WIDTH_RANGE

//---------------------------------------------------------------------------------------------------------------------
// NoC (external) Ports Information

`define NOC_CONT_NOC_NUM_OF_PORTS          4

`define NOC_CONT_NOC_NUM_OF_PORTS_VECTOR_RANGE       `NOC_CONT_NOC_NUM_OF_PORTS-1 : 0
`define NOC_CONT_NOC_NUM_OF_PKT_DEST_VECTOR_RANGE    `NOC_CONT_NOC_NUM_OF_PORTS : 0    // destinations are local plus ports 0-3

`define NOC_CONT_NOC_NUM_OF_PORTS_MSB     (`CLOG2(`NOC_CONT_NOC_NUM_OF_PORTS))
`define NOC_CONT_NOC_NUM_OF_PORTS_LSB     0
`define NOC_CONT_NOC_NUM_OF_PORTS_SIZE    (`NOC_CONT_NOC_NUM_OF_PORTS_MSB - `NOC_CONT_NOC_NUM_OF_PORTS_LSB +1)
`define NOC_CONT_NOC_NUM_OF_PORTS_RANGE    `NOC_CONT_NOC_NUM_OF_PORTS_MSB : `NOC_CONT_NOC_NUM_OF_PORTS_LSB

`define NOC_CONT_NOC_PROTOCOL_CNTL_SOP            1
`define NOC_CONT_NOC_PROTOCOL_CNTL_DATA           0
`define NOC_CONT_NOC_PROTOCOL_CNTL_EOP            2
`define NOC_CONT_NOC_PROTOCOL_CNTL_SOP_EOP        3

`define NOC_CONT_NOC_PROTOCOL_CNTL_SOD            1
`define NOC_CONT_NOC_PROTOCOL_CNTL_EOD            2
`define NOC_CONT_NOC_PROTOCOL_CNTL_SOD_EOD        3

// Port signalling
`define NOC_CONT_NOC_PORT_CNTL_WIDTH               2
`define NOC_CONT_NOC_PORT_CNTL_MSB                 `NOC_CONT_NOC_PORT_CNTL_WIDTH-1
`define NOC_CONT_NOC_PORT_CNTL_LSB                 0
`define NOC_CONT_NOC_PORT_CNTL_RANGE               `NOC_CONT_NOC_PORT_CNTL_MSB : `NOC_CONT_NOC_PORT_CNTL_LSB

`define NOC_CONT_NOC_PORT_DATA_WIDTH               `NOC_CONT_EXTERNAL_DATA_WIDTH         
`define NOC_CONT_NOC_PORT_DATA_MSB                 `NOC_CONT_NOC_PORT_DATA_WIDTH-1
`define NOC_CONT_NOC_PORT_DATA_LSB                 0
`define NOC_CONT_NOC_PORT_DATA_RANGE               `NOC_CONT_NOC_PORT_DATA_MSB : `NOC_CONT_NOC_PORT_DATA_LSB



//---------------------------------------------------------------------------------------------------------------------
//---------------------------------------------------------------------------------------------------------------------
// FSM(s) 

// Local Input Queue Controller
`include "/home/lbbaker/Cortical/StreamingOps/PE/HDL/common/noc_cntl_noc_local_inq_control_fsm_state_definitions.vh"

// Local Output Queue Controller
`define NOC_CONT_LOCAL_OUTQ_CNTL_WAIT                    15'b000_0000_0000_0001
`define NOC_CONT_LOCAL_OUTQ_CNTL_CP_FIFO_READ            15'b000_0000_0000_0010
`define NOC_CONT_LOCAL_OUTQ_CNTL_CP_PORT_REQ             15'b000_0000_0000_0100
`define NOC_CONT_LOCAL_OUTQ_CNTL_CP_SEND_HEADER          15'b000_0000_0000_1000
`define NOC_CONT_LOCAL_OUTQ_CNTL_CP_SEND_CYCLE2          15'b000_0000_0001_0000
`define NOC_CONT_LOCAL_OUTQ_CNTL_CP_SEND_CYCLE3          15'b000_0000_0010_0000
`define NOC_CONT_LOCAL_OUTQ_CNTL_CP_COMPLETE             15'b000_0000_0100_0000
`define NOC_CONT_LOCAL_OUTQ_CNTL_DP_FIFO_READ            15'b000_0000_1000_0000
`define NOC_CONT_LOCAL_OUTQ_CNTL_DP_PORT_REQ             15'b000_0001_0000_0000
`define NOC_CONT_LOCAL_OUTQ_CNTL_DP_SEND_HEADER          15'b000_0010_0000_0000
`define NOC_CONT_LOCAL_OUTQ_CNTL_DP_SEND_CYCLE2          15'b000_0100_0000_0000
`define NOC_CONT_LOCAL_OUTQ_CNTL_DP_SEND_CYCLE3          15'b000_1000_0000_0000
`define NOC_CONT_LOCAL_OUTQ_CNTL_DP_COMPLETE             15'b001_0000_0000_0000
`define NOC_CONT_LOCAL_OUTQ_CNTL_COMPLETE                15'b010_0000_0000_0000
`define NOC_CONT_LOCAL_OUTQ_CNTL_ERROR                   15'b100_0000_0000_0000

`define NOC_CONT_LOCAL_OUTQ_CNTL_STATE_MSB          14
`define NOC_CONT_LOCAL_OUTQ_CNTL_STATE_LSB           0
`define NOC_CONT_LOCAL_OUTQ_CNTL_STATE_SIZE          (`NOC_CONT_LOCAL_OUTQ_CNTL_STATE_MSB - `NOC_CONT_LOCAL_OUTQ_CNTL_STATE_LSB +1)
`define NOC_CONT_LOCAL_OUTQ_CNTL_STATE_RANGE          `NOC_CONT_LOCAL_OUTQ_CNTL_STATE_MSB : `NOC_CONT_LOCAL_OUTQ_CNTL_STATE_LSB


// Port Output Controller
`include "/home/lbbaker/Cortical/StreamingOps/PE/HDL/common/noc_cntl_noc_port_output_control_fsm_state_definitions.vh"


// Port Input Controller
`define NOC_CONT_NOC_PORT_INPUT_CNTL_WAIT                     7'b000_0001
`define NOC_CONT_NOC_PORT_INPUT_CNTL_FIFO_READ                7'b000_0010
`define NOC_CONT_NOC_PORT_INPUT_CNTL_DESTINATION_REQ          7'b000_0100
`define NOC_CONT_NOC_PORT_INPUT_CNTL_TRANSFER_HEADER          7'b000_1000
`define NOC_CONT_NOC_PORT_INPUT_CNTL_TRANSFER_PACKET          7'b001_0000
`define NOC_CONT_NOC_PORT_INPUT_CNTL_COMPLETE                 7'b010_0000
`define NOC_CONT_NOC_PORT_INPUT_CNTL_ERROR                    7'b100_0000

`define NOC_CONT_NOC_PORT_INPUT_CNTL_STATE_MSB           6
`define NOC_CONT_NOC_PORT_INPUT_CNTL_STATE_LSB           0
`define NOC_CONT_NOC_PORT_INPUT_CNTL_STATE_SIZE          (`NOC_CONT_NOC_PORT_INPUT_CNTL_STATE_MSB - `NOC_CONT_NOC_PORT_INPUT_CNTL_STATE_LSB +1)
`define NOC_CONT_NOC_PORT_INPUT_CNTL_STATE_RANGE          `NOC_CONT_NOC_PORT_INPUT_CNTL_STATE_MSB : `NOC_CONT_NOC_PORT_INPUT_CNTL_STATE_LSB


// end of FSM(s)
//---------------------------------------------------------------------------------------------------------------------
//---------------------------------------------------------------------------------------------------------------------

//---------------------------------------------------------------------------------------------------------------------
//---------------------------------------------------------------------------------------------------------------------
// Packet Types

`define NOC_CONT_TYPE_STATUS            0
`define NOC_CONT_TYPE_WRITE_REQUEST     1
`define NOC_CONT_TYPE_DMA_REQUEST       2
`define NOC_CONT_TYPE_READ_REQUEST      3
`define NOC_CONT_TYPE_READ_RESPONCE     4
`define NOC_CONT_TYPE_DMA_DATA          5
`define NOC_CONT_TYPE_DMA_DATA_SOD      6
`define NOC_CONT_TYPE_DMA_DATA_EOD      7

// Destination address types

`define NOC_CONT_DESTINATION_ADDR_TYPE_BITMASK           0
`define NOC_CONT_DESTINATION_ADDR_TYPE_MCAST_GROUP       1
`define NOC_CONT_DESTINATION_ADDR_TYPE_UNICAST           2

//---------------------------------------------------------------------------------------------------------------------
// First Cycle of all NoC packets are the same (external fields)

// 1st Transaction on external bus
`define NOC_CONT_EXTERNAL_1ST_CYCLE_PAD_SIZE                1
`define NOC_CONT_EXTERNAL_1ST_CYCLE_PAD_MSB                 `NOC_CONT_EXTERNAL_1ST_CYCLE_PAD_SIZE-1
`define NOC_CONT_EXTERNAL_1ST_CYCLE_PAD_LSB                 0
`define NOC_CONT_EXTERNAL_1ST_CYCLE_PAD_RANGE               `NOC_CONT_EXTERNAL_1ST_CYCLE_PAD_MSB : `NOC_CONT_EXTERNAL_1ST_CYCLE_PAD_LSB

`define NOC_CONT_EXTERNAL_1ST_CYCLE_PRIORITY_SIZE                1
`define NOC_CONT_EXTERNAL_1ST_CYCLE_PRIORITY_MSB                 (`NOC_CONT_EXTERNAL_1ST_CYCLE_PRIORITY_LSB + `NOC_CONT_EXTERNAL_1ST_CYCLE_PRIORITY_SIZE-1)
`define NOC_CONT_EXTERNAL_1ST_CYCLE_PRIORITY_LSB                 (`NOC_CONT_EXTERNAL_1ST_CYCLE_PAD_MSB + 1)
`define NOC_CONT_EXTERNAL_1ST_CYCLE_PRIORITY_RANGE               `NOC_CONT_EXTERNAL_1ST_CYCLE_PRIORITY_MSB : `NOC_CONT_EXTERNAL_1ST_CYCLE_PRIORITY_LSB
`define NOC_CONT_EXTERNAL_1ST_CYCLE_PRIORITY_CP              0
`define NOC_CONT_EXTERNAL_1ST_CYCLE_PRIORITY_DP              1

`define NOC_CONT_EXTERNAL_1ST_CYCLE_DESTINATION_ADDR_SIZE                 32
`define NOC_CONT_EXTERNAL_1ST_CYCLE_DESTINATION_ADDR_MSB                   (`NOC_CONT_EXTERNAL_1ST_CYCLE_DESTINATION_ADDR_LSB + `NOC_CONT_EXTERNAL_1ST_CYCLE_DESTINATION_ADDR_SIZE-1)
`define NOC_CONT_EXTERNAL_1ST_CYCLE_DESTINATION_ADDR_LSB                   (`NOC_CONT_EXTERNAL_1ST_CYCLE_PRIORITY_MSB + 1)
`define NOC_CONT_EXTERNAL_1ST_CYCLE_DESTINATION_ADDR_RANGE                 `NOC_CONT_EXTERNAL_1ST_CYCLE_DESTINATION_ADDR_MSB : `NOC_CONT_EXTERNAL_1ST_CYCLE_DESTINATION_ADDR_LSB

`define NOC_CONT_EXTERNAL_1ST_CYCLE_DESTINATION_ADDR_TYPE_SIZE                  2
`define NOC_CONT_EXTERNAL_1ST_CYCLE_DESTINATION_ADDR_TYPE_MSB                   (`NOC_CONT_EXTERNAL_1ST_CYCLE_DESTINATION_ADDR_TYPE_LSB + `NOC_CONT_EXTERNAL_1ST_CYCLE_DESTINATION_ADDR_TYPE_SIZE-1)
`define NOC_CONT_EXTERNAL_1ST_CYCLE_DESTINATION_ADDR_TYPE_LSB                   (`NOC_CONT_EXTERNAL_1ST_CYCLE_DESTINATION_ADDR_MSB + 1)
`define NOC_CONT_EXTERNAL_1ST_CYCLE_DESTINATION_ADDR_TYPE_RANGE                 `NOC_CONT_EXTERNAL_1ST_CYCLE_DESTINATION_ADDR_TYPE_MSB : `NOC_CONT_EXTERNAL_1ST_CYCLE_DESTINATION_ADDR_TYPE_LSB

`define NOC_CONT_EXTERNAL_1ST_CYCLE_SOURCE_PE_SIZE                  6
`define NOC_CONT_EXTERNAL_1ST_CYCLE_SOURCE_PE_MSB                   (`NOC_CONT_EXTERNAL_1ST_CYCLE_SOURCE_PE_LSB + `NOC_CONT_EXTERNAL_1ST_CYCLE_SOURCE_PE_SIZE-1)
`define NOC_CONT_EXTERNAL_1ST_CYCLE_SOURCE_PE_LSB                   (`NOC_CONT_EXTERNAL_1ST_CYCLE_DESTINATION_ADDR_TYPE_MSB + 1)
`define NOC_CONT_EXTERNAL_1ST_CYCLE_SOURCE_PE_RANGE                 `NOC_CONT_EXTERNAL_1ST_CYCLE_SOURCE_PE_MSB : `NOC_CONT_EXTERNAL_1ST_CYCLE_SOURCE_PE_LSB


//---------------------------------------------------------------------------------------------------------------------
// DMA Request (external fields)

// Fields
`define NOC_CONT_NOC_PACKET_TYPE_MSB            3
`define NOC_CONT_NOC_PACKET_TYPE_LSB            0
`define NOC_CONT_NOC_PACKET_TYPE_SIZE           (`NOC_CONT_NOC_PACKET_TYPE_MSB - `NOC_CONT_NOC_PACKET_TYPE_LSB +1)
`define NOC_CONT_NOC_PACKET_TYPE_RANGE           `NOC_CONT_NOC_PACKET_TYPE_MSB : `NOC_CONT_NOC_PACKET_TYPE_LSB

`define NOC_CONT_EXTERNAL_DMA_WORDS_PER_PKT                16

// 2nd Transaction on external bus
`define NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_PAD_SIZE                1
`define NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_PAD_MSB                 `NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_PAD_SIZE-1
`define NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_PAD_LSB                 0
`define NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_PAD_RANGE               `NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_PAD_MSB : `NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_PAD_LSB

`define NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_STAGGER_SIZE                  8
`define NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_STAGGER_MSB                   (`NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_STAGGER_LSB + `NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_STAGGER_SIZE-1)
`define NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_STAGGER_LSB                   (`NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_PAD_MSB + 1)
`define NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_STAGGER_RANGE                 `NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_STAGGER_MSB : `NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_STAGGER_LSB

`define NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_ADDRESS_SIZE                 24
`define NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_ADDRESS_MSB                   (`NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_ADDRESS_LSB + `NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_ADDRESS_SIZE-1)
`define NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_ADDRESS_LSB                   (`NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_STAGGER_MSB + 1)
`define NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_ADDRESS_RANGE                 `NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_ADDRESS_MSB : `NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_ADDRESS_LSB

`define NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_STRM_ID_SIZE                  1
`define NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_STRM_ID_MSB                   (`NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_STRM_ID_LSB + `NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_STRM_ID_SIZE-1)
`define NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_STRM_ID_LSB                   (`NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_ADDRESS_MSB + 1)
`define NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_STRM_ID_RANGE                 `NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_STRM_ID_MSB : `NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_STRM_ID_LSB

`define NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_LANE_ID_SIZE                  4
`define NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_LANE_ID_MSB                   (`NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_LANE_ID_LSB + `NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_LANE_ID_SIZE-1)
`define NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_LANE_ID_LSB                   (`NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_STRM_ID_MSB + 1)
`define NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_LANE_ID_RANGE                 `NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_LANE_ID_MSB : `NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_LANE_ID_LSB

`define NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_TYPE_SIZE                  4
`define NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_TYPE_MSB                   (`NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_TYPE_LSB + `NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_TYPE_SIZE-1)
`define NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_TYPE_LSB                   (`NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_LANE_ID_MSB + 1)
`define NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_TYPE_RANGE                 `NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_TYPE_MSB : `NOC_CONT_EXTERNAL_DMA_REQ_2ND_CYCLE_TYPE_LSB

// 3rd Transaction on external bus
`define NOC_CONT_EXTERNAL_DMA_REQ_3RD_CYCLE_PAD_SIZE                18
`define NOC_CONT_EXTERNAL_DMA_REQ_3RD_CYCLE_PAD_MSB                 `NOC_CONT_EXTERNAL_DMA_REQ_3RD_CYCLE_PAD_SIZE-1
`define NOC_CONT_EXTERNAL_DMA_REQ_3RD_CYCLE_PAD_LSB                 0
`define NOC_CONT_EXTERNAL_DMA_REQ_3RD_CYCLE_PAD_RANGE               `NOC_CONT_EXTERNAL_DMA_REQ_3RD_CYCLE_PAD_MSB : `NOC_CONT_EXTERNAL_DMA_REQ_3RD_CYCLE_PAD_LSB

`define NOC_CONT_EXTERNAL_DMA_REQ_3RD_CYCLE_NUM_OF_WORDS_SIZE             20
`define NOC_CONT_EXTERNAL_DMA_REQ_3RD_CYCLE_NUM_OF_WORDS_MSB              (`NOC_CONT_EXTERNAL_DMA_REQ_3RD_CYCLE_NUM_OF_WORDS_LSB + `NOC_CONT_EXTERNAL_DMA_REQ_3RD_CYCLE_NUM_OF_WORDS_SIZE-1)
`define NOC_CONT_EXTERNAL_DMA_REQ_3RD_CYCLE_NUM_OF_WORDS_LSB              (`NOC_CONT_EXTERNAL_DMA_REQ_3RD_CYCLE_PAD_MSB + 1)
`define NOC_CONT_EXTERNAL_DMA_REQ_3RD_CYCLE_NUM_OF_WORDS_RANGE            `NOC_CONT_EXTERNAL_DMA_REQ_3RD_CYCLE_NUM_OF_WORDS_MSB : `NOC_CONT_EXTERNAL_DMA_REQ_3RD_CYCLE_NUM_OF_WORDS_LSB

`define NOC_CONT_EXTERNAL_DMA_REQ_3RD_CYCLE_PAYLOAD_TYPE_SIZE             4
`define NOC_CONT_EXTERNAL_DMA_REQ_3RD_CYCLE_PAYLOAD_TYPE_MSB              (`NOC_CONT_EXTERNAL_DMA_REQ_3RD_CYCLE_PAYLOAD_TYPE_LSB + `NOC_CONT_EXTERNAL_DMA_REQ_3RD_CYCLE_PAYLOAD_TYPE_SIZE-1)
`define NOC_CONT_EXTERNAL_DMA_REQ_3RD_CYCLE_PAYLOAD_TYPE_LSB              (`NOC_CONT_EXTERNAL_DMA_REQ_3RD_CYCLE_NUM_OF_WORDS_MSB + 1)
`define NOC_CONT_EXTERNAL_DMA_REQ_3RD_CYCLE_PAYLOAD_TYPE_RANGE            `NOC_CONT_EXTERNAL_DMA_REQ_3RD_CYCLE_PAYLOAD_TYPE_MSB : `NOC_CONT_EXTERNAL_DMA_REQ_3RD_CYCLE_PAYLOAD_TYPE_LSB

//---------------------------------------------------------------------------------------------------------------------
// DMA Request (internal fields)

`define NOC_CONT_INTERNAL_DMA_WORDS_PER_PKT                16

// First Transaction on internal bus
`define NOC_CONT_INTERNAL_DMA_REQ_1ST_CYCLE_PAD_SIZE                8
`define NOC_CONT_INTERNAL_DMA_REQ_1ST_CYCLE_PAD_MSB                 `NOC_CONT_INTERNAL_DMA_REQ_1ST_CYCLE_PAD_SIZE-1
`define NOC_CONT_INTERNAL_DMA_REQ_1ST_CYCLE_PAD_LSB                 0
`define NOC_CONT_INTERNAL_DMA_REQ_1ST_CYCLE_PAD_RANGE               `NOC_CONT_INTERNAL_DMA_REQ_1ST_CYCLE_PAD_MSB : `NOC_CONT_INTERNAL_DMA_REQ_1ST_CYCLE_PAD_LSB

`define NOC_CONT_INTERNAL_DMA_REQ_1ST_CYCLE_STAGGER_SIZE                  8
`define NOC_CONT_INTERNAL_DMA_REQ_1ST_CYCLE_STAGGER_MSB                   (`NOC_CONT_INTERNAL_DMA_REQ_1ST_CYCLE_STAGGER_LSB + `NOC_CONT_INTERNAL_DMA_REQ_1ST_CYCLE_STAGGER_SIZE-1)
`define NOC_CONT_INTERNAL_DMA_REQ_1ST_CYCLE_STAGGER_LSB                   (`NOC_CONT_INTERNAL_DMA_REQ_1ST_CYCLE_PAD_MSB + 1)
`define NOC_CONT_INTERNAL_DMA_REQ_1ST_CYCLE_STAGGER_RANGE                 `NOC_CONT_INTERNAL_DMA_REQ_1ST_CYCLE_STAGGER_MSB : `NOC_CONT_INTERNAL_DMA_REQ_1ST_CYCLE_STAGGER_LSB

`define NOC_CONT_INTERNAL_DMA_REQ_1ST_CYCLE_ADDRESS_SIZE                 24
`define NOC_CONT_INTERNAL_DMA_REQ_1ST_CYCLE_ADDRESS_MSB                   (`NOC_CONT_INTERNAL_DMA_REQ_1ST_CYCLE_ADDRESS_LSB + `NOC_CONT_INTERNAL_DMA_REQ_1ST_CYCLE_ADDRESS_SIZE-1)
`define NOC_CONT_INTERNAL_DMA_REQ_1ST_CYCLE_ADDRESS_LSB                   (`NOC_CONT_INTERNAL_DMA_REQ_1ST_CYCLE_STAGGER_MSB + 1)
`define NOC_CONT_INTERNAL_DMA_REQ_1ST_CYCLE_ADDRESS_RANGE                 `NOC_CONT_INTERNAL_DMA_REQ_1ST_CYCLE_ADDRESS_MSB : `NOC_CONT_INTERNAL_DMA_REQ_1ST_CYCLE_ADDRESS_LSB

// Second Transaction on internal bus
`define NOC_CONT_INTERNAL_DMA_REQ_2ND_CYCLE_PAD_SIZE                16
`define NOC_CONT_INTERNAL_DMA_REQ_2ND_CYCLE_PAD_MSB                 `NOC_CONT_INTERNAL_DMA_REQ_2ND_CYCLE_PAD_SIZE-1
`define NOC_CONT_INTERNAL_DMA_REQ_2ND_CYCLE_PAD_LSB                 0
`define NOC_CONT_INTERNAL_DMA_REQ_2ND_CYCLE_PAD_RANGE               `NOC_CONT_INTERNAL_DMA_REQ_2ND_CYCLE_PAD_MSB : `NOC_CONT_INTERNAL_DMA_REQ_2ND_CYCLE_PAD_LSB

`define NOC_CONT_INTERNAL_DMA_REQ_2ND_CYCLE_NUM_OF_WORDS_SIZE             20
`define NOC_CONT_INTERNAL_DMA_REQ_2ND_CYCLE_NUM_OF_WORDS_MSB              (`NOC_CONT_INTERNAL_DMA_REQ_2ND_CYCLE_NUM_OF_WORDS_LSB + `NOC_CONT_INTERNAL_DMA_REQ_2ND_CYCLE_NUM_OF_WORDS_SIZE-1)
`define NOC_CONT_INTERNAL_DMA_REQ_2ND_CYCLE_NUM_OF_WORDS_LSB              (`NOC_CONT_INTERNAL_DMA_REQ_2ND_CYCLE_PAD_MSB + 1)
`define NOC_CONT_INTERNAL_DMA_REQ_2ND_CYCLE_NUM_OF_WORDS_RANGE            `NOC_CONT_INTERNAL_DMA_REQ_2ND_CYCLE_NUM_OF_WORDS_MSB : `NOC_CONT_INTERNAL_DMA_REQ_2ND_CYCLE_NUM_OF_WORDS_LSB

`define NOC_CONT_INTERNAL_DMA_REQ_2ND_CYCLE_PAYLOAD_TYPE_SIZE             4
`define NOC_CONT_INTERNAL_DMA_REQ_2ND_CYCLE_PAYLOAD_TYPE_MSB              (`NOC_CONT_INTERNAL_DMA_REQ_2ND_CYCLE_PAYLOAD_TYPE_LSB + `NOC_CONT_INTERNAL_DMA_REQ_2ND_CYCLE_PAYLOAD_TYPE_SIZE-1)
`define NOC_CONT_INTERNAL_DMA_REQ_2ND_CYCLE_PAYLOAD_TYPE_LSB              (`NOC_CONT_INTERNAL_DMA_REQ_2ND_CYCLE_NUM_OF_WORDS_MSB + 1)
`define NOC_CONT_INTERNAL_DMA_REQ_2ND_CYCLE_PAYLOAD_TYPE_RANGE            `NOC_CONT_INTERNAL_DMA_REQ_2ND_CYCLE_PAYLOAD_TYPE_MSB : `NOC_CONT_INTERNAL_DMA_REQ_2ND_CYCLE_PAYLOAD_TYPE_LSB


//---------------------------------------------------------------------------------------------------------------------
// DMA Data (external fields)

// First transactions on internal bus
`define NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_DATA_SIZE                32
`define NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_DATA_MSB                 `NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_DATA_SIZE-1
`define NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_DATA_LSB                 0
`define NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_DATA_RANGE               `NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_DATA_MSB : `NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_DATA_LSB

`define NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_4OR8_SIZE                  1
`define NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_4OR8_MSB                   (`NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_4OR8_LSB + `NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_4OR8_SIZE-1)
`define NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_4OR8_LSB                   (`NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_DATA_MSB + 1)
`define NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_4OR8_RANGE                 `NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_4OR8_MSB : `NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_4OR8_LSB

`define NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_STRM_ID_SIZE                  1
`define NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_STRM_ID_MSB                   (`NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_STRM_ID_LSB + `NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_STRM_ID_SIZE-1)
`define NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_STRM_ID_LSB                   (`NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_4OR8_MSB + 1)
`define NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_STRM_ID_RANGE                 `NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_STRM_ID_MSB : `NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_STRM_ID_LSB

`define NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_LANE_ID_SIZE                  4
`define NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_LANE_ID_MSB                   (`NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_LANE_ID_LSB + `NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_LANE_ID_SIZE-1)
`define NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_LANE_ID_LSB                   (`NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_STRM_ID_MSB + 1)
`define NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_LANE_ID_RANGE                 `NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_LANE_ID_MSB : `NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_LANE_ID_LSB

`define NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_TYPE_SIZE                  4
`define NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_TYPE_MSB                   (`NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_TYPE_LSB + `NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_TYPE_SIZE-1)
`define NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_TYPE_LSB                   (`NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_LANE_ID_MSB + 1)
`define NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_TYPE_RANGE                 `NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_TYPE_MSB : `NOC_CONT_EXTERNAL_DMA_DATA_2ND_CYCLE_TYPE_LSB

// All other transactions on internal bus
`define NOC_CONT_EXTERNAL_DMA_DATA_ALL_CYCLE_DATA_SIZE                32
`define NOC_CONT_EXTERNAL_DMA_DATA_ALL_CYCLE_DATA_MSB                 `NOC_CONT_EXTERNAL_DMA_DATA_ALL_CYCLE_DATA_SIZE-1
`define NOC_CONT_EXTERNAL_DMA_DATA_ALL_CYCLE_DATA_LSB                 0
`define NOC_CONT_EXTERNAL_DMA_DATA_ALL_CYCLE_DATA_RANGE               `NOC_CONT_EXTERNAL_DMA_DATA_ALL_CYCLE_DATA_MSB : `NOC_CONT_EXTERNAL_DMA_DATA_ALL_CYCLE_DATA_LSB

`define NOC_CONT_EXTERNAL_DMA_DATA_ALL_CYCLE_PAD_SIZE                  10
`define NOC_CONT_EXTERNAL_DMA_DATA_ALL_CYCLE_PAD_MSB                   (`NOC_CONT_EXTERNAL_DMA_DATA_ALL_CYCLE_PAD_LSB + `NOC_CONT_EXTERNAL_DMA_DATA_ALL_CYCLE_PAD_SIZE-1)
`define NOC_CONT_EXTERNAL_DMA_DATA_ALL_CYCLE_PAD_LSB                   (`NOC_CONT_EXTERNAL_DMA_DATA_ALL_CYCLE_DATA_MSB + 1)
`define NOC_CONT_EXTERNAL_DMA_DATA_ALL_CYCLE_PAD_RANGE                 `NOC_CONT_EXTERNAL_DMA_DATA_ALL_CYCLE_PAD_MSB : `NOC_CONT_EXTERNAL_DMA_DATA_ALL_CYCLE_PAD_LSB


//---------------------------------------------------------------------------------------------------------------------
// DMA Data (internal fields)

// First transactions on internal bus
`define NOC_CONT_INTERNAL_DMA_DATA_1ST_CYCLE_DATA_SIZE                32
`define NOC_CONT_INTERNAL_DMA_DATA_1ST_CYCLE_DATA_MSB                 `NOC_CONT_INTERNAL_DMA_DATA_1ST_CYCLE_DATA_SIZE-1
`define NOC_CONT_INTERNAL_DMA_DATA_1ST_CYCLE_DATA_LSB                 0
`define NOC_CONT_INTERNAL_DMA_DATA_1ST_CYCLE_DATA_RANGE               `NOC_CONT_INTERNAL_DMA_DATA_1ST_CYCLE_DATA_MSB : `NOC_CONT_INTERNAL_DMA_DATA_1ST_CYCLE_DATA_LSB

`define NOC_CONT_INTERNAL_DMA_DATA_1ST_CYCLE_4OR8_SIZE                  1
`define NOC_CONT_INTERNAL_DMA_DATA_1ST_CYCLE_4OR8_MSB                   (`NOC_CONT_INTERNAL_DMA_DATA_1ST_CYCLE_4OR8_LSB + `NOC_CONT_INTERNAL_DMA_DATA_1ST_CYCLE_4OR8_SIZE-1)
`define NOC_CONT_INTERNAL_DMA_DATA_1ST_CYCLE_4OR8_LSB                   (`NOC_CONT_INTERNAL_DMA_DATA_1ST_CYCLE_DATA_MSB + 1)
`define NOC_CONT_INTERNAL_DMA_DATA_1ST_CYCLE_4OR8_RANGE                 `NOC_CONT_INTERNAL_DMA_DATA_1ST_CYCLE_4OR8_MSB : `NOC_CONT_INTERNAL_DMA_DATA_1ST_CYCLE_4OR8_LSB

`define NOC_CONT_INTERNAL_DMA_DATA_1ST_CYCLE_PAD_SIZE                  7
`define NOC_CONT_INTERNAL_DMA_DATA_1ST_CYCLE_PAD_MSB                   (`NOC_CONT_INTERNAL_DMA_DATA_1ST_CYCLE_PAD_LSB + `NOC_CONT_INTERNAL_DMA_DATA_1ST_CYCLE_PAD_SIZE-1)
`define NOC_CONT_INTERNAL_DMA_DATA_1ST_CYCLE_PAD_LSB                   (`NOC_CONT_INTERNAL_DMA_DATA_1ST_CYCLE_4OR8_MSB + 1)
`define NOC_CONT_INTERNAL_DMA_DATA_1ST_CYCLE_PAD_RANGE                 `NOC_CONT_INTERNAL_DMA_DATA_1ST_CYCLE_PAD_MSB : `NOC_CONT_INTERNAL_DMA_DATA_1ST_CYCLE_PAD_LSB

// All other transactions on internal bus
`define NOC_CONT_INTERNAL_DMA_DATA_ALL_CYCLE_DATA_SIZE                32
`define NOC_CONT_INTERNAL_DMA_DATA_ALL_CYCLE_DATA_MSB                 `NOC_CONT_INTERNAL_DMA_DATA_ALL_CYCLE_DATA_SIZE-1
`define NOC_CONT_INTERNAL_DMA_DATA_ALL_CYCLE_DATA_LSB                 0
`define NOC_CONT_INTERNAL_DMA_DATA_ALL_CYCLE_DATA_RANGE               `NOC_CONT_INTERNAL_DMA_DATA_ALL_CYCLE_DATA_MSB : `NOC_CONT_INTERNAL_DMA_DATA_ALL_CYCLE_DATA_LSB

`define NOC_CONT_INTERNAL_DMA_DATA_ALL_CYCLE_PAD_SIZE                  8
`define NOC_CONT_INTERNAL_DMA_DATA_ALL_CYCLE_PAD_MSB                   (`NOC_CONT_INTERNAL_DMA_DATA_ALL_CYCLE_PAD_LSB + `NOC_CONT_INTERNAL_DMA_DATA_ALL_CYCLE_PAD_SIZE-1)
`define NOC_CONT_INTERNAL_DMA_DATA_ALL_CYCLE_PAD_LSB                   (`NOC_CONT_INTERNAL_DMA_DATA_ALL_CYCLE_DATA_MSB + 1)
`define NOC_CONT_INTERNAL_DMA_DATA_ALL_CYCLE_PAD_RANGE                 `NOC_CONT_INTERNAL_DMA_DATA_ALL_CYCLE_PAD_MSB : `NOC_CONT_INTERNAL_DMA_DATA_ALL_CYCLE_PAD_LSB


// end of Packet Types
//---------------------------------------------------------------------------------------------------------------------
//---------------------------------------------------------------------------------------------------------------------

//------------------------------------------------
// Internal to NoC Interface data FIFO
//------------------------------------------------

`define NOC_CONT_TO_INTF_DATA_FIFO_DEPTH          32
`define NOC_CONT_TO_INTF_DATA_FIFO_DEPTH_MSB      (`NOC_CONT_TO_INTF_DATA_FIFO_DEPTH) -1
`define NOC_CONT_TO_INTF_DATA_FIFO_DEPTH_LSB      0
`define NOC_CONT_TO_INTF_DATA_FIFO_DEPTH_SIZE     (`NOC_CONT_TO_INTF_DATA_FIFO_DEPTH_MSB - `NOC_CONT_TO_INTF_DATA_FIFO_DEPTH_LSB +1)
`define NOC_CONT_TO_INTF_DATA_FIFO_DEPTH_RANGE     `NOC_CONT_TO_INTF_DATA_FIFO_DEPTH_MSB : `NOC_CONT_TO_INTF_DATA_FIFO_DEPTH_LSB
`define NOC_CONT_TO_INTF_DATA_FIFO_MSB            ((`CLOG2(`NOC_CONT_TO_INTF_DATA_FIFO_DEPTH)) -1)
`define NOC_CONT_TO_INTF_DATA_FIFO_LSB            0
`define NOC_CONT_TO_INTF_DATA_FIFO_SIZE           (`NOC_CONT_TO_INTF_DATA_FIFO_MSB - `NOC_CONT_TO_INTF_DATA_FIFO_LSB +1)
`define NOC_CONT_TO_INTF_DATA_FIFO_RANGE           `NOC_CONT_TO_INTF_DATA_FIFO_MSB : `NOC_CONT_TO_INTF_DATA_FIFO_LSB

// Count number of packets in internal datapath FIFO
`define NOC_CONT_TO_INTF_DATA_FIFO_EOP_COUNT_MSB     2
`define NOC_CONT_TO_INTF_DATA_FIFO_EOP_COUNT_LSB     0
`define NOC_CONT_TO_INTF_DATA_FIFO_EOP_COUNT_SIZE    (`NOC_CONT_TO_INTF_DATA_FIFO_EOP_COUNT_MSB - `NOC_CONT_TO_INTF_DATA_FIFO_EOP_COUNT_LSB +1)
`define NOC_CONT_TO_INTF_DATA_FIFO_EOP_COUNT_RANGE    `NOC_CONT_TO_INTF_DATA_FIFO_EOP_COUNT_MSB : `NOC_CONT_TO_INTF_DATA_FIFO_EOP_COUNT_LSB

//------------------------------------------------
// External from NoC Interface Control FIFO
//------------------------------------------------

`define NOC_CONT_FROM_EXT_NOC_CNTL_FIFO_DEPTH          64
`define NOC_CONT_FROM_EXT_NOC_CNTL_FIFO_DEPTH_MSB      (`NOC_CONT_FROM_EXT_NOC_CNTL_FIFO_DEPTH) -1
`define NOC_CONT_FROM_EXT_NOC_CNTL_FIFO_DEPTH_LSB      0
`define NOC_CONT_FROM_EXT_NOC_CNTL_FIFO_DEPTH_SIZE     (`NOC_CONT_FROM_EXT_NOC_CNTL_FIFO_DEPTH_MSB - `NOC_CONT_FROM_EXT_NOC_CNTL_FIFO_DEPTH_LSB +1)
`define NOC_CONT_FROM_EXT_NOC_CNTL_FIFO_DEPTH_RANGE     `NOC_CONT_FROM_EXT_NOC_CNTL_FIFO_DEPTH_MSB : `NOC_CONT_FROM_EXT_NOC_CNTL_FIFO_DEPTH_LSB
`define NOC_CONT_FROM_EXT_NOC_CNTL_FIFO_MSB            ((`CLOG2(`NOC_CONT_FROM_EXT_NOC_CNTL_FIFO_DEPTH)) -1)
`define NOC_CONT_FROM_EXT_NOC_CNTL_FIFO_LSB            0
`define NOC_CONT_FROM_EXT_NOC_CNTL_FIFO_SIZE           (`NOC_CONT_FROM_EXT_NOC_CNTL_FIFO_MSB - `NOC_CONT_FROM_EXT_NOC_CNTL_FIFO_LSB +1)
`define NOC_CONT_FROM_EXT_NOC_CNTL_FIFO_RANGE           `NOC_CONT_FROM_EXT_NOC_CNTL_FIFO_MSB : `NOC_CONT_FROM_EXT_NOC_CNTL_FIFO_LSB

// Threshold below full when we assert almost full
`define NOC_CONT_FROM_EXT_NOC_CNTL_FIFO_ALMOST_FULL_THRESHOLD  6

// Count number of packets in internal datapath FIFO
`define NOC_CONT_FROM_EXT_NOC_CNTL_FIFO_EOP_COUNT_MSB     8
`define NOC_CONT_FROM_EXT_NOC_CNTL_FIFO_EOP_COUNT_LSB     0
`define NOC_CONT_FROM_EXT_NOC_CNTL_FIFO_EOP_COUNT_SIZE    (`NOC_CONT_FROM_EXT_NOC_CNTL_FIFO_EOP_COUNT_MSB - `NOC_CONT_FROM_EXT_NOC_CNTL_FIFO_EOP_COUNT_LSB +1)
`define NOC_CONT_FROM_EXT_NOC_CNTL_FIFO_EOP_COUNT_RANGE    `NOC_CONT_FROM_EXT_NOC_CNTL_FIFO_EOP_COUNT_MSB : `NOC_CONT_FROM_EXT_NOC_CNTL_FIFO_EOP_COUNT_LSB

