
            // Common (Scalar) Register(s)                
            .simd__cntl__rs0         ( simd__cntl__rs0        ),
            .simd__cntl__rs1         ( simd__cntl__rs1        ),

            // Lane 31             
            .simd__cntl__lane_r128   ( simd__cntl__lane_r128  ),
            .simd__cntl__lane_r129   ( simd__cntl__lane_r129  ),
            .simd__cntl__lane_r130   ( simd__cntl__lane_r130  ),
            .simd__cntl__lane_r131   ( simd__cntl__lane_r131  ),
            .simd__cntl__lane_r132   ( simd__cntl__lane_r132  ),
            .simd__cntl__lane_r133   ( simd__cntl__lane_r133  ),
            .simd__cntl__lane_r134   ( simd__cntl__lane_r134  ),
            .simd__cntl__lane_r135   ( simd__cntl__lane_r135  ),
