
            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe0__oob_cntl                         ( std__pe0__oob_cntl   ),
            .std__pe0__oob_valid                        ( std__pe0__oob_valid  ),
            .pe0__std__oob_ready                        ( pe0__std__oob_ready  ),
            .std__pe0__oob_type                         ( std__pe0__oob_type   ),
            .std__pe0__oob_data                         ( std__pe0__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe1__oob_cntl                         ( std__pe1__oob_cntl   ),
            .std__pe1__oob_valid                        ( std__pe1__oob_valid  ),
            .pe1__std__oob_ready                        ( pe1__std__oob_ready  ),
            .std__pe1__oob_type                         ( std__pe1__oob_type   ),
            .std__pe1__oob_data                         ( std__pe1__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe2__oob_cntl                         ( std__pe2__oob_cntl   ),
            .std__pe2__oob_valid                        ( std__pe2__oob_valid  ),
            .pe2__std__oob_ready                        ( pe2__std__oob_ready  ),
            .std__pe2__oob_type                         ( std__pe2__oob_type   ),
            .std__pe2__oob_data                         ( std__pe2__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe3__oob_cntl                         ( std__pe3__oob_cntl   ),
            .std__pe3__oob_valid                        ( std__pe3__oob_valid  ),
            .pe3__std__oob_ready                        ( pe3__std__oob_ready  ),
            .std__pe3__oob_type                         ( std__pe3__oob_type   ),
            .std__pe3__oob_data                         ( std__pe3__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe4__oob_cntl                         ( std__pe4__oob_cntl   ),
            .std__pe4__oob_valid                        ( std__pe4__oob_valid  ),
            .pe4__std__oob_ready                        ( pe4__std__oob_ready  ),
            .std__pe4__oob_type                         ( std__pe4__oob_type   ),
            .std__pe4__oob_data                         ( std__pe4__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe5__oob_cntl                         ( std__pe5__oob_cntl   ),
            .std__pe5__oob_valid                        ( std__pe5__oob_valid  ),
            .pe5__std__oob_ready                        ( pe5__std__oob_ready  ),
            .std__pe5__oob_type                         ( std__pe5__oob_type   ),
            .std__pe5__oob_data                         ( std__pe5__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe6__oob_cntl                         ( std__pe6__oob_cntl   ),
            .std__pe6__oob_valid                        ( std__pe6__oob_valid  ),
            .pe6__std__oob_ready                        ( pe6__std__oob_ready  ),
            .std__pe6__oob_type                         ( std__pe6__oob_type   ),
            .std__pe6__oob_data                         ( std__pe6__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe7__oob_cntl                         ( std__pe7__oob_cntl   ),
            .std__pe7__oob_valid                        ( std__pe7__oob_valid  ),
            .pe7__std__oob_ready                        ( pe7__std__oob_ready  ),
            .std__pe7__oob_type                         ( std__pe7__oob_type   ),
            .std__pe7__oob_data                         ( std__pe7__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe8__oob_cntl                         ( std__pe8__oob_cntl   ),
            .std__pe8__oob_valid                        ( std__pe8__oob_valid  ),
            .pe8__std__oob_ready                        ( pe8__std__oob_ready  ),
            .std__pe8__oob_type                         ( std__pe8__oob_type   ),
            .std__pe8__oob_data                         ( std__pe8__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe9__oob_cntl                         ( std__pe9__oob_cntl   ),
            .std__pe9__oob_valid                        ( std__pe9__oob_valid  ),
            .pe9__std__oob_ready                        ( pe9__std__oob_ready  ),
            .std__pe9__oob_type                         ( std__pe9__oob_type   ),
            .std__pe9__oob_data                         ( std__pe9__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe10__oob_cntl                         ( std__pe10__oob_cntl   ),
            .std__pe10__oob_valid                        ( std__pe10__oob_valid  ),
            .pe10__std__oob_ready                        ( pe10__std__oob_ready  ),
            .std__pe10__oob_type                         ( std__pe10__oob_type   ),
            .std__pe10__oob_data                         ( std__pe10__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe11__oob_cntl                         ( std__pe11__oob_cntl   ),
            .std__pe11__oob_valid                        ( std__pe11__oob_valid  ),
            .pe11__std__oob_ready                        ( pe11__std__oob_ready  ),
            .std__pe11__oob_type                         ( std__pe11__oob_type   ),
            .std__pe11__oob_data                         ( std__pe11__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe12__oob_cntl                         ( std__pe12__oob_cntl   ),
            .std__pe12__oob_valid                        ( std__pe12__oob_valid  ),
            .pe12__std__oob_ready                        ( pe12__std__oob_ready  ),
            .std__pe12__oob_type                         ( std__pe12__oob_type   ),
            .std__pe12__oob_data                         ( std__pe12__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe13__oob_cntl                         ( std__pe13__oob_cntl   ),
            .std__pe13__oob_valid                        ( std__pe13__oob_valid  ),
            .pe13__std__oob_ready                        ( pe13__std__oob_ready  ),
            .std__pe13__oob_type                         ( std__pe13__oob_type   ),
            .std__pe13__oob_data                         ( std__pe13__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe14__oob_cntl                         ( std__pe14__oob_cntl   ),
            .std__pe14__oob_valid                        ( std__pe14__oob_valid  ),
            .pe14__std__oob_ready                        ( pe14__std__oob_ready  ),
            .std__pe14__oob_type                         ( std__pe14__oob_type   ),
            .std__pe14__oob_data                         ( std__pe14__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe15__oob_cntl                         ( std__pe15__oob_cntl   ),
            .std__pe15__oob_valid                        ( std__pe15__oob_valid  ),
            .pe15__std__oob_ready                        ( pe15__std__oob_ready  ),
            .std__pe15__oob_type                         ( std__pe15__oob_type   ),
            .std__pe15__oob_data                         ( std__pe15__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe16__oob_cntl                         ( std__pe16__oob_cntl   ),
            .std__pe16__oob_valid                        ( std__pe16__oob_valid  ),
            .pe16__std__oob_ready                        ( pe16__std__oob_ready  ),
            .std__pe16__oob_type                         ( std__pe16__oob_type   ),
            .std__pe16__oob_data                         ( std__pe16__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe17__oob_cntl                         ( std__pe17__oob_cntl   ),
            .std__pe17__oob_valid                        ( std__pe17__oob_valid  ),
            .pe17__std__oob_ready                        ( pe17__std__oob_ready  ),
            .std__pe17__oob_type                         ( std__pe17__oob_type   ),
            .std__pe17__oob_data                         ( std__pe17__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe18__oob_cntl                         ( std__pe18__oob_cntl   ),
            .std__pe18__oob_valid                        ( std__pe18__oob_valid  ),
            .pe18__std__oob_ready                        ( pe18__std__oob_ready  ),
            .std__pe18__oob_type                         ( std__pe18__oob_type   ),
            .std__pe18__oob_data                         ( std__pe18__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe19__oob_cntl                         ( std__pe19__oob_cntl   ),
            .std__pe19__oob_valid                        ( std__pe19__oob_valid  ),
            .pe19__std__oob_ready                        ( pe19__std__oob_ready  ),
            .std__pe19__oob_type                         ( std__pe19__oob_type   ),
            .std__pe19__oob_data                         ( std__pe19__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe20__oob_cntl                         ( std__pe20__oob_cntl   ),
            .std__pe20__oob_valid                        ( std__pe20__oob_valid  ),
            .pe20__std__oob_ready                        ( pe20__std__oob_ready  ),
            .std__pe20__oob_type                         ( std__pe20__oob_type   ),
            .std__pe20__oob_data                         ( std__pe20__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe21__oob_cntl                         ( std__pe21__oob_cntl   ),
            .std__pe21__oob_valid                        ( std__pe21__oob_valid  ),
            .pe21__std__oob_ready                        ( pe21__std__oob_ready  ),
            .std__pe21__oob_type                         ( std__pe21__oob_type   ),
            .std__pe21__oob_data                         ( std__pe21__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe22__oob_cntl                         ( std__pe22__oob_cntl   ),
            .std__pe22__oob_valid                        ( std__pe22__oob_valid  ),
            .pe22__std__oob_ready                        ( pe22__std__oob_ready  ),
            .std__pe22__oob_type                         ( std__pe22__oob_type   ),
            .std__pe22__oob_data                         ( std__pe22__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe23__oob_cntl                         ( std__pe23__oob_cntl   ),
            .std__pe23__oob_valid                        ( std__pe23__oob_valid  ),
            .pe23__std__oob_ready                        ( pe23__std__oob_ready  ),
            .std__pe23__oob_type                         ( std__pe23__oob_type   ),
            .std__pe23__oob_data                         ( std__pe23__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe24__oob_cntl                         ( std__pe24__oob_cntl   ),
            .std__pe24__oob_valid                        ( std__pe24__oob_valid  ),
            .pe24__std__oob_ready                        ( pe24__std__oob_ready  ),
            .std__pe24__oob_type                         ( std__pe24__oob_type   ),
            .std__pe24__oob_data                         ( std__pe24__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe25__oob_cntl                         ( std__pe25__oob_cntl   ),
            .std__pe25__oob_valid                        ( std__pe25__oob_valid  ),
            .pe25__std__oob_ready                        ( pe25__std__oob_ready  ),
            .std__pe25__oob_type                         ( std__pe25__oob_type   ),
            .std__pe25__oob_data                         ( std__pe25__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe26__oob_cntl                         ( std__pe26__oob_cntl   ),
            .std__pe26__oob_valid                        ( std__pe26__oob_valid  ),
            .pe26__std__oob_ready                        ( pe26__std__oob_ready  ),
            .std__pe26__oob_type                         ( std__pe26__oob_type   ),
            .std__pe26__oob_data                         ( std__pe26__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe27__oob_cntl                         ( std__pe27__oob_cntl   ),
            .std__pe27__oob_valid                        ( std__pe27__oob_valid  ),
            .pe27__std__oob_ready                        ( pe27__std__oob_ready  ),
            .std__pe27__oob_type                         ( std__pe27__oob_type   ),
            .std__pe27__oob_data                         ( std__pe27__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe28__oob_cntl                         ( std__pe28__oob_cntl   ),
            .std__pe28__oob_valid                        ( std__pe28__oob_valid  ),
            .pe28__std__oob_ready                        ( pe28__std__oob_ready  ),
            .std__pe28__oob_type                         ( std__pe28__oob_type   ),
            .std__pe28__oob_data                         ( std__pe28__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe29__oob_cntl                         ( std__pe29__oob_cntl   ),
            .std__pe29__oob_valid                        ( std__pe29__oob_valid  ),
            .pe29__std__oob_ready                        ( pe29__std__oob_ready  ),
            .std__pe29__oob_type                         ( std__pe29__oob_type   ),
            .std__pe29__oob_data                         ( std__pe29__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe30__oob_cntl                         ( std__pe30__oob_cntl   ),
            .std__pe30__oob_valid                        ( std__pe30__oob_valid  ),
            .pe30__std__oob_ready                        ( pe30__std__oob_ready  ),
            .std__pe30__oob_type                         ( std__pe30__oob_type   ),
            .std__pe30__oob_data                         ( std__pe30__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe31__oob_cntl                         ( std__pe31__oob_cntl   ),
            .std__pe31__oob_valid                        ( std__pe31__oob_valid  ),
            .pe31__std__oob_ready                        ( pe31__std__oob_ready  ),
            .std__pe31__oob_type                         ( std__pe31__oob_type   ),
            .std__pe31__oob_data                         ( std__pe31__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe32__oob_cntl                         ( std__pe32__oob_cntl   ),
            .std__pe32__oob_valid                        ( std__pe32__oob_valid  ),
            .pe32__std__oob_ready                        ( pe32__std__oob_ready  ),
            .std__pe32__oob_type                         ( std__pe32__oob_type   ),
            .std__pe32__oob_data                         ( std__pe32__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe33__oob_cntl                         ( std__pe33__oob_cntl   ),
            .std__pe33__oob_valid                        ( std__pe33__oob_valid  ),
            .pe33__std__oob_ready                        ( pe33__std__oob_ready  ),
            .std__pe33__oob_type                         ( std__pe33__oob_type   ),
            .std__pe33__oob_data                         ( std__pe33__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe34__oob_cntl                         ( std__pe34__oob_cntl   ),
            .std__pe34__oob_valid                        ( std__pe34__oob_valid  ),
            .pe34__std__oob_ready                        ( pe34__std__oob_ready  ),
            .std__pe34__oob_type                         ( std__pe34__oob_type   ),
            .std__pe34__oob_data                         ( std__pe34__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe35__oob_cntl                         ( std__pe35__oob_cntl   ),
            .std__pe35__oob_valid                        ( std__pe35__oob_valid  ),
            .pe35__std__oob_ready                        ( pe35__std__oob_ready  ),
            .std__pe35__oob_type                         ( std__pe35__oob_type   ),
            .std__pe35__oob_data                         ( std__pe35__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe36__oob_cntl                         ( std__pe36__oob_cntl   ),
            .std__pe36__oob_valid                        ( std__pe36__oob_valid  ),
            .pe36__std__oob_ready                        ( pe36__std__oob_ready  ),
            .std__pe36__oob_type                         ( std__pe36__oob_type   ),
            .std__pe36__oob_data                         ( std__pe36__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe37__oob_cntl                         ( std__pe37__oob_cntl   ),
            .std__pe37__oob_valid                        ( std__pe37__oob_valid  ),
            .pe37__std__oob_ready                        ( pe37__std__oob_ready  ),
            .std__pe37__oob_type                         ( std__pe37__oob_type   ),
            .std__pe37__oob_data                         ( std__pe37__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe38__oob_cntl                         ( std__pe38__oob_cntl   ),
            .std__pe38__oob_valid                        ( std__pe38__oob_valid  ),
            .pe38__std__oob_ready                        ( pe38__std__oob_ready  ),
            .std__pe38__oob_type                         ( std__pe38__oob_type   ),
            .std__pe38__oob_data                         ( std__pe38__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe39__oob_cntl                         ( std__pe39__oob_cntl   ),
            .std__pe39__oob_valid                        ( std__pe39__oob_valid  ),
            .pe39__std__oob_ready                        ( pe39__std__oob_ready  ),
            .std__pe39__oob_type                         ( std__pe39__oob_type   ),
            .std__pe39__oob_data                         ( std__pe39__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe40__oob_cntl                         ( std__pe40__oob_cntl   ),
            .std__pe40__oob_valid                        ( std__pe40__oob_valid  ),
            .pe40__std__oob_ready                        ( pe40__std__oob_ready  ),
            .std__pe40__oob_type                         ( std__pe40__oob_type   ),
            .std__pe40__oob_data                         ( std__pe40__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe41__oob_cntl                         ( std__pe41__oob_cntl   ),
            .std__pe41__oob_valid                        ( std__pe41__oob_valid  ),
            .pe41__std__oob_ready                        ( pe41__std__oob_ready  ),
            .std__pe41__oob_type                         ( std__pe41__oob_type   ),
            .std__pe41__oob_data                         ( std__pe41__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe42__oob_cntl                         ( std__pe42__oob_cntl   ),
            .std__pe42__oob_valid                        ( std__pe42__oob_valid  ),
            .pe42__std__oob_ready                        ( pe42__std__oob_ready  ),
            .std__pe42__oob_type                         ( std__pe42__oob_type   ),
            .std__pe42__oob_data                         ( std__pe42__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe43__oob_cntl                         ( std__pe43__oob_cntl   ),
            .std__pe43__oob_valid                        ( std__pe43__oob_valid  ),
            .pe43__std__oob_ready                        ( pe43__std__oob_ready  ),
            .std__pe43__oob_type                         ( std__pe43__oob_type   ),
            .std__pe43__oob_data                         ( std__pe43__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe44__oob_cntl                         ( std__pe44__oob_cntl   ),
            .std__pe44__oob_valid                        ( std__pe44__oob_valid  ),
            .pe44__std__oob_ready                        ( pe44__std__oob_ready  ),
            .std__pe44__oob_type                         ( std__pe44__oob_type   ),
            .std__pe44__oob_data                         ( std__pe44__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe45__oob_cntl                         ( std__pe45__oob_cntl   ),
            .std__pe45__oob_valid                        ( std__pe45__oob_valid  ),
            .pe45__std__oob_ready                        ( pe45__std__oob_ready  ),
            .std__pe45__oob_type                         ( std__pe45__oob_type   ),
            .std__pe45__oob_data                         ( std__pe45__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe46__oob_cntl                         ( std__pe46__oob_cntl   ),
            .std__pe46__oob_valid                        ( std__pe46__oob_valid  ),
            .pe46__std__oob_ready                        ( pe46__std__oob_ready  ),
            .std__pe46__oob_type                         ( std__pe46__oob_type   ),
            .std__pe46__oob_data                         ( std__pe46__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe47__oob_cntl                         ( std__pe47__oob_cntl   ),
            .std__pe47__oob_valid                        ( std__pe47__oob_valid  ),
            .pe47__std__oob_ready                        ( pe47__std__oob_ready  ),
            .std__pe47__oob_type                         ( std__pe47__oob_type   ),
            .std__pe47__oob_data                         ( std__pe47__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe48__oob_cntl                         ( std__pe48__oob_cntl   ),
            .std__pe48__oob_valid                        ( std__pe48__oob_valid  ),
            .pe48__std__oob_ready                        ( pe48__std__oob_ready  ),
            .std__pe48__oob_type                         ( std__pe48__oob_type   ),
            .std__pe48__oob_data                         ( std__pe48__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe49__oob_cntl                         ( std__pe49__oob_cntl   ),
            .std__pe49__oob_valid                        ( std__pe49__oob_valid  ),
            .pe49__std__oob_ready                        ( pe49__std__oob_ready  ),
            .std__pe49__oob_type                         ( std__pe49__oob_type   ),
            .std__pe49__oob_data                         ( std__pe49__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe50__oob_cntl                         ( std__pe50__oob_cntl   ),
            .std__pe50__oob_valid                        ( std__pe50__oob_valid  ),
            .pe50__std__oob_ready                        ( pe50__std__oob_ready  ),
            .std__pe50__oob_type                         ( std__pe50__oob_type   ),
            .std__pe50__oob_data                         ( std__pe50__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe51__oob_cntl                         ( std__pe51__oob_cntl   ),
            .std__pe51__oob_valid                        ( std__pe51__oob_valid  ),
            .pe51__std__oob_ready                        ( pe51__std__oob_ready  ),
            .std__pe51__oob_type                         ( std__pe51__oob_type   ),
            .std__pe51__oob_data                         ( std__pe51__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe52__oob_cntl                         ( std__pe52__oob_cntl   ),
            .std__pe52__oob_valid                        ( std__pe52__oob_valid  ),
            .pe52__std__oob_ready                        ( pe52__std__oob_ready  ),
            .std__pe52__oob_type                         ( std__pe52__oob_type   ),
            .std__pe52__oob_data                         ( std__pe52__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe53__oob_cntl                         ( std__pe53__oob_cntl   ),
            .std__pe53__oob_valid                        ( std__pe53__oob_valid  ),
            .pe53__std__oob_ready                        ( pe53__std__oob_ready  ),
            .std__pe53__oob_type                         ( std__pe53__oob_type   ),
            .std__pe53__oob_data                         ( std__pe53__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe54__oob_cntl                         ( std__pe54__oob_cntl   ),
            .std__pe54__oob_valid                        ( std__pe54__oob_valid  ),
            .pe54__std__oob_ready                        ( pe54__std__oob_ready  ),
            .std__pe54__oob_type                         ( std__pe54__oob_type   ),
            .std__pe54__oob_data                         ( std__pe54__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe55__oob_cntl                         ( std__pe55__oob_cntl   ),
            .std__pe55__oob_valid                        ( std__pe55__oob_valid  ),
            .pe55__std__oob_ready                        ( pe55__std__oob_ready  ),
            .std__pe55__oob_type                         ( std__pe55__oob_type   ),
            .std__pe55__oob_data                         ( std__pe55__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe56__oob_cntl                         ( std__pe56__oob_cntl   ),
            .std__pe56__oob_valid                        ( std__pe56__oob_valid  ),
            .pe56__std__oob_ready                        ( pe56__std__oob_ready  ),
            .std__pe56__oob_type                         ( std__pe56__oob_type   ),
            .std__pe56__oob_data                         ( std__pe56__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe57__oob_cntl                         ( std__pe57__oob_cntl   ),
            .std__pe57__oob_valid                        ( std__pe57__oob_valid  ),
            .pe57__std__oob_ready                        ( pe57__std__oob_ready  ),
            .std__pe57__oob_type                         ( std__pe57__oob_type   ),
            .std__pe57__oob_data                         ( std__pe57__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe58__oob_cntl                         ( std__pe58__oob_cntl   ),
            .std__pe58__oob_valid                        ( std__pe58__oob_valid  ),
            .pe58__std__oob_ready                        ( pe58__std__oob_ready  ),
            .std__pe58__oob_type                         ( std__pe58__oob_type   ),
            .std__pe58__oob_data                         ( std__pe58__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe59__oob_cntl                         ( std__pe59__oob_cntl   ),
            .std__pe59__oob_valid                        ( std__pe59__oob_valid  ),
            .pe59__std__oob_ready                        ( pe59__std__oob_ready  ),
            .std__pe59__oob_type                         ( std__pe59__oob_type   ),
            .std__pe59__oob_data                         ( std__pe59__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe60__oob_cntl                         ( std__pe60__oob_cntl   ),
            .std__pe60__oob_valid                        ( std__pe60__oob_valid  ),
            .pe60__std__oob_ready                        ( pe60__std__oob_ready  ),
            .std__pe60__oob_type                         ( std__pe60__oob_type   ),
            .std__pe60__oob_data                         ( std__pe60__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe61__oob_cntl                         ( std__pe61__oob_cntl   ),
            .std__pe61__oob_valid                        ( std__pe61__oob_valid  ),
            .pe61__std__oob_ready                        ( pe61__std__oob_ready  ),
            .std__pe61__oob_type                         ( std__pe61__oob_type   ),
            .std__pe61__oob_data                         ( std__pe61__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe62__oob_cntl                         ( std__pe62__oob_cntl   ),
            .std__pe62__oob_valid                        ( std__pe62__oob_valid  ),
            .pe62__std__oob_ready                        ( pe62__std__oob_ready  ),
            .std__pe62__oob_type                         ( std__pe62__oob_type   ),
            .std__pe62__oob_data                         ( std__pe62__oob_data   ),


            // OOB controls the PE                         
            // For now assume OOB is separate to lanes     
            .std__pe63__oob_cntl                         ( std__pe63__oob_cntl   ),
            .std__pe63__oob_valid                        ( std__pe63__oob_valid  ),
            .pe63__std__oob_ready                        ( pe63__std__oob_ready  ),
            .std__pe63__oob_type                         ( std__pe63__oob_type   ),
            .std__pe63__oob_data                         ( std__pe63__oob_data   ),

