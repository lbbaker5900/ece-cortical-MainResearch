
        wire                                      read_data_strm_valid_next  ;  
        reg                                       read_data_strm_valid       ;  