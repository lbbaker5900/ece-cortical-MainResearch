
            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr0__std__oob_cntl                         ( mgr0__std__oob_cntl   ),
            .mgr0__std__oob_valid                        ( mgr0__std__oob_valid  ),
            .std__mgr0__oob_ready                        ( std__mgr0__oob_ready  ),
            .mgr0__std__oob_type                         ( mgr0__std__oob_type   ),
            .mgr0__std__oob_data                         ( mgr0__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr1__std__oob_cntl                         ( mgr1__std__oob_cntl   ),
            .mgr1__std__oob_valid                        ( mgr1__std__oob_valid  ),
            .std__mgr1__oob_ready                        ( std__mgr1__oob_ready  ),
            .mgr1__std__oob_type                         ( mgr1__std__oob_type   ),
            .mgr1__std__oob_data                         ( mgr1__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr2__std__oob_cntl                         ( mgr2__std__oob_cntl   ),
            .mgr2__std__oob_valid                        ( mgr2__std__oob_valid  ),
            .std__mgr2__oob_ready                        ( std__mgr2__oob_ready  ),
            .mgr2__std__oob_type                         ( mgr2__std__oob_type   ),
            .mgr2__std__oob_data                         ( mgr2__std__oob_data   ),

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            .mgr3__std__oob_cntl                         ( mgr3__std__oob_cntl   ),
            .mgr3__std__oob_valid                        ( mgr3__std__oob_valid  ),
            .std__mgr3__oob_ready                        ( std__mgr3__oob_ready  ),
            .mgr3__std__oob_type                         ( mgr3__std__oob_type   ),
            .mgr3__std__oob_data                         ( mgr3__std__oob_data   ),
