
    force pe_array_inst.pe_inst[0].pe.simd__scntl__rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r128 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r129 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r130 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r131 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[0].pe.ldst__memc__request        = 1'b0 ; 
    force pe_array_inst.pe_inst[0].pe.ldst__memc__released       = 1'b1 ; 
    force pe_array_inst.pe_inst[0].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[0].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[0].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[0].pe.ldst__memc__write_valid    = 1'b0; 
    force pe_array_inst.pe_inst[0].pe.ldst__memc__read_valid     = 1'b0; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r128 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r129 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r130 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r131 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[1].pe.ldst__memc__request        = 1'b0 ; 
    force pe_array_inst.pe_inst[1].pe.ldst__memc__released       = 1'b1 ; 
    force pe_array_inst.pe_inst[1].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[1].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[1].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[1].pe.ldst__memc__write_valid    = 1'b0; 
    force pe_array_inst.pe_inst[1].pe.ldst__memc__read_valid     = 1'b0; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r128 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r129 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r130 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r131 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[2].pe.ldst__memc__request        = 1'b0 ; 
    force pe_array_inst.pe_inst[2].pe.ldst__memc__released       = 1'b1 ; 
    force pe_array_inst.pe_inst[2].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[2].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[2].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[2].pe.ldst__memc__write_valid    = 1'b0; 
    force pe_array_inst.pe_inst[2].pe.ldst__memc__read_valid     = 1'b0; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__rs0        = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__rs1        = 32'b1111_1111_1111_1111_1111_1111_1111_1111; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [0] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [1] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [2] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [3] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [4] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [5] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [6] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [7] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [8] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [9] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [10] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [11] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [12] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [13] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [14] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [15] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [16] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [17] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [18] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [19] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [20] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [21] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [22] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [23] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [24] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [25] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [26] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [27] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [28] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [29] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [30] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r128 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r129 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r130 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r131 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [31] = 32'b0000_0000_0000_0000_0000_0000_0000_0000; 
    force pe_array_inst.pe_inst[3].pe.ldst__memc__request        = 1'b0 ; 
    force pe_array_inst.pe_inst[3].pe.ldst__memc__released       = 1'b1 ; 
    force pe_array_inst.pe_inst[3].pe.ldst__memc__write_address  = 'd0 ; 
    force pe_array_inst.pe_inst[3].pe.ldst__memc__write_data     = 'd0 ; 
    force pe_array_inst.pe_inst[3].pe.ldst__memc__read_address   = 'h00 ; 
    force pe_array_inst.pe_inst[3].pe.ldst__memc__write_valid    = 1'b0; 
    force pe_array_inst.pe_inst[3].pe.ldst__memc__read_valid     = 1'b0; 