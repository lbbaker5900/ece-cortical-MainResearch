
  // NoC port 0
  .mgr__noc__port0_valid           ( mgr__noc__port0_valid           ),
  .mgr__noc__port0_cntl            ( mgr__noc__port0_cntl            ),
  .mgr__noc__port0_data            ( mgr__noc__port0_data            ),
  .noc__mgr__port0_fc              ( noc__mgr__port0_fc              ),
  .noc__mgr__port0_valid           ( noc__mgr__port0_valid           ),
  .noc__mgr__port0_cntl            ( noc__mgr__port0_cntl            ),
  .noc__mgr__port0_data            ( noc__mgr__port0_data            ),
  .mgr__noc__port0_fc              ( mgr__noc__port0_fc              ),
  .sys__mgr__port0_destinationMask ( sys__mgr__port0_destinationMask ),

  // NoC port 1
  .mgr__noc__port1_valid           ( mgr__noc__port1_valid           ),
  .mgr__noc__port1_cntl            ( mgr__noc__port1_cntl            ),
  .mgr__noc__port1_data            ( mgr__noc__port1_data            ),
  .noc__mgr__port1_fc              ( noc__mgr__port1_fc              ),
  .noc__mgr__port1_valid           ( noc__mgr__port1_valid           ),
  .noc__mgr__port1_cntl            ( noc__mgr__port1_cntl            ),
  .noc__mgr__port1_data            ( noc__mgr__port1_data            ),
  .mgr__noc__port1_fc              ( mgr__noc__port1_fc              ),
  .sys__mgr__port1_destinationMask ( sys__mgr__port1_destinationMask ),

  // NoC port 2
  .mgr__noc__port2_valid           ( mgr__noc__port2_valid           ),
  .mgr__noc__port2_cntl            ( mgr__noc__port2_cntl            ),
  .mgr__noc__port2_data            ( mgr__noc__port2_data            ),
  .noc__mgr__port2_fc              ( noc__mgr__port2_fc              ),
  .noc__mgr__port2_valid           ( noc__mgr__port2_valid           ),
  .noc__mgr__port2_cntl            ( noc__mgr__port2_cntl            ),
  .noc__mgr__port2_data            ( noc__mgr__port2_data            ),
  .mgr__noc__port2_fc              ( mgr__noc__port2_fc              ),
  .sys__mgr__port2_destinationMask ( sys__mgr__port2_destinationMask ),

  // NoC port 3
  .mgr__noc__port3_valid           ( mgr__noc__port3_valid           ),
  .mgr__noc__port3_cntl            ( mgr__noc__port3_cntl            ),
  .mgr__noc__port3_data            ( mgr__noc__port3_data            ),
  .noc__mgr__port3_fc              ( noc__mgr__port3_fc              ),
  .noc__mgr__port3_valid           ( noc__mgr__port3_valid           ),
  .noc__mgr__port3_cntl            ( noc__mgr__port3_cntl            ),
  .noc__mgr__port3_data            ( noc__mgr__port3_data            ),
  .mgr__noc__port3_fc              ( mgr__noc__port3_fc              ),
  .sys__mgr__port3_destinationMask ( sys__mgr__port3_destinationMask ),

