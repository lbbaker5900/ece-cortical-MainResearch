
    1 :  // note: in system verilog checker, we increment cycle count 1..8 not 0..7
      begin
        upstream_packet_data [0] = upstream_data[31:0] ; 
        upstream_packet_data [1] = upstream_data[63:32] ; 
        upstream_packet_data [2] = upstream_data[95:64] ; 
        upstream_packet_data [3] = upstream_data[127:96] ; 
      end 
    2 :  // note: in system verilog checker, we increment cycle count 1..8 not 0..7
      begin
        upstream_packet_data [4] = upstream_data[31:0] ; 
        upstream_packet_data [5] = upstream_data[63:32] ; 
        upstream_packet_data [6] = upstream_data[95:64] ; 
        upstream_packet_data [7] = upstream_data[127:96] ; 
      end 
    3 :  // note: in system verilog checker, we increment cycle count 1..8 not 0..7
      begin
        upstream_packet_data [8] = upstream_data[31:0] ; 
        upstream_packet_data [9] = upstream_data[63:32] ; 
        upstream_packet_data [10] = upstream_data[95:64] ; 
        upstream_packet_data [11] = upstream_data[127:96] ; 
      end 
    4 :  // note: in system verilog checker, we increment cycle count 1..8 not 0..7
      begin
        upstream_packet_data [12] = upstream_data[31:0] ; 
        upstream_packet_data [13] = upstream_data[63:32] ; 
        upstream_packet_data [14] = upstream_data[95:64] ; 
        upstream_packet_data [15] = upstream_data[127:96] ; 
      end 
    5 :  // note: in system verilog checker, we increment cycle count 1..8 not 0..7
      begin
        upstream_packet_data [16] = upstream_data[31:0] ; 
        upstream_packet_data [17] = upstream_data[63:32] ; 
        upstream_packet_data [18] = upstream_data[95:64] ; 
        upstream_packet_data [19] = upstream_data[127:96] ; 
      end 
    6 :  // note: in system verilog checker, we increment cycle count 1..8 not 0..7
      begin
        upstream_packet_data [20] = upstream_data[31:0] ; 
        upstream_packet_data [21] = upstream_data[63:32] ; 
        upstream_packet_data [22] = upstream_data[95:64] ; 
        upstream_packet_data [23] = upstream_data[127:96] ; 
      end 
    7 :  // note: in system verilog checker, we increment cycle count 1..8 not 0..7
      begin
        upstream_packet_data [24] = upstream_data[31:0] ; 
        upstream_packet_data [25] = upstream_data[63:32] ; 
        upstream_packet_data [26] = upstream_data[95:64] ; 
        upstream_packet_data [27] = upstream_data[127:96] ; 
      end 
    8 :  // note: in system verilog checker, we increment cycle count 1..8 not 0..7
      begin
        upstream_packet_data [28] = upstream_data[31:0] ; 
        upstream_packet_data [29] = upstream_data[63:32] ; 
        upstream_packet_data [30] = upstream_data[95:64] ; 
        upstream_packet_data [31] = upstream_data[127:96] ; 
      end 