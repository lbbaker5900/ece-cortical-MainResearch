
    .reg__scntl__lane0_ready   ( reg__scntl__lane0_ready  ) ,
    .scntl__reg__lane0_valid   ( scntl__reg__lane0_valid  ) ,
    .scntl__reg__lane0_cntl    ( scntl__reg__lane0_cntl   ) ,
    .scntl__reg__lane0_data    ( scntl__reg__lane0_data   ) ,

    .reg__scntl__lane1_ready   ( reg__scntl__lane1_ready  ) ,
    .scntl__reg__lane1_valid   ( scntl__reg__lane1_valid  ) ,
    .scntl__reg__lane1_cntl    ( scntl__reg__lane1_cntl   ) ,
    .scntl__reg__lane1_data    ( scntl__reg__lane1_data   ) ,

    .reg__scntl__lane2_ready   ( reg__scntl__lane2_ready  ) ,
    .scntl__reg__lane2_valid   ( scntl__reg__lane2_valid  ) ,
    .scntl__reg__lane2_cntl    ( scntl__reg__lane2_cntl   ) ,
    .scntl__reg__lane2_data    ( scntl__reg__lane2_data   ) ,

    .reg__scntl__lane3_ready   ( reg__scntl__lane3_ready  ) ,
    .scntl__reg__lane3_valid   ( scntl__reg__lane3_valid  ) ,
    .scntl__reg__lane3_cntl    ( scntl__reg__lane3_cntl   ) ,
    .scntl__reg__lane3_data    ( scntl__reg__lane3_data   ) ,

    .reg__scntl__lane4_ready   ( reg__scntl__lane4_ready  ) ,
    .scntl__reg__lane4_valid   ( scntl__reg__lane4_valid  ) ,
    .scntl__reg__lane4_cntl    ( scntl__reg__lane4_cntl   ) ,
    .scntl__reg__lane4_data    ( scntl__reg__lane4_data   ) ,

    .reg__scntl__lane5_ready   ( reg__scntl__lane5_ready  ) ,
    .scntl__reg__lane5_valid   ( scntl__reg__lane5_valid  ) ,
    .scntl__reg__lane5_cntl    ( scntl__reg__lane5_cntl   ) ,
    .scntl__reg__lane5_data    ( scntl__reg__lane5_data   ) ,

    .reg__scntl__lane6_ready   ( reg__scntl__lane6_ready  ) ,
    .scntl__reg__lane6_valid   ( scntl__reg__lane6_valid  ) ,
    .scntl__reg__lane6_cntl    ( scntl__reg__lane6_cntl   ) ,
    .scntl__reg__lane6_data    ( scntl__reg__lane6_data   ) ,

    .reg__scntl__lane7_ready   ( reg__scntl__lane7_ready  ) ,
    .scntl__reg__lane7_valid   ( scntl__reg__lane7_valid  ) ,
    .scntl__reg__lane7_cntl    ( scntl__reg__lane7_cntl   ) ,
    .scntl__reg__lane7_data    ( scntl__reg__lane7_data   ) ,

    .reg__scntl__lane8_ready   ( reg__scntl__lane8_ready  ) ,
    .scntl__reg__lane8_valid   ( scntl__reg__lane8_valid  ) ,
    .scntl__reg__lane8_cntl    ( scntl__reg__lane8_cntl   ) ,
    .scntl__reg__lane8_data    ( scntl__reg__lane8_data   ) ,

    .reg__scntl__lane9_ready   ( reg__scntl__lane9_ready  ) ,
    .scntl__reg__lane9_valid   ( scntl__reg__lane9_valid  ) ,
    .scntl__reg__lane9_cntl    ( scntl__reg__lane9_cntl   ) ,
    .scntl__reg__lane9_data    ( scntl__reg__lane9_data   ) ,

    .reg__scntl__lane10_ready   ( reg__scntl__lane10_ready  ) ,
    .scntl__reg__lane10_valid   ( scntl__reg__lane10_valid  ) ,
    .scntl__reg__lane10_cntl    ( scntl__reg__lane10_cntl   ) ,
    .scntl__reg__lane10_data    ( scntl__reg__lane10_data   ) ,

    .reg__scntl__lane11_ready   ( reg__scntl__lane11_ready  ) ,
    .scntl__reg__lane11_valid   ( scntl__reg__lane11_valid  ) ,
    .scntl__reg__lane11_cntl    ( scntl__reg__lane11_cntl   ) ,
    .scntl__reg__lane11_data    ( scntl__reg__lane11_data   ) ,

    .reg__scntl__lane12_ready   ( reg__scntl__lane12_ready  ) ,
    .scntl__reg__lane12_valid   ( scntl__reg__lane12_valid  ) ,
    .scntl__reg__lane12_cntl    ( scntl__reg__lane12_cntl   ) ,
    .scntl__reg__lane12_data    ( scntl__reg__lane12_data   ) ,

    .reg__scntl__lane13_ready   ( reg__scntl__lane13_ready  ) ,
    .scntl__reg__lane13_valid   ( scntl__reg__lane13_valid  ) ,
    .scntl__reg__lane13_cntl    ( scntl__reg__lane13_cntl   ) ,
    .scntl__reg__lane13_data    ( scntl__reg__lane13_data   ) ,

    .reg__scntl__lane14_ready   ( reg__scntl__lane14_ready  ) ,
    .scntl__reg__lane14_valid   ( scntl__reg__lane14_valid  ) ,
    .scntl__reg__lane14_cntl    ( scntl__reg__lane14_cntl   ) ,
    .scntl__reg__lane14_data    ( scntl__reg__lane14_data   ) ,

    .reg__scntl__lane15_ready   ( reg__scntl__lane15_ready  ) ,
    .scntl__reg__lane15_valid   ( scntl__reg__lane15_valid  ) ,
    .scntl__reg__lane15_cntl    ( scntl__reg__lane15_cntl   ) ,
    .scntl__reg__lane15_data    ( scntl__reg__lane15_data   ) ,

    .reg__scntl__lane16_ready   ( reg__scntl__lane16_ready  ) ,
    .scntl__reg__lane16_valid   ( scntl__reg__lane16_valid  ) ,
    .scntl__reg__lane16_cntl    ( scntl__reg__lane16_cntl   ) ,
    .scntl__reg__lane16_data    ( scntl__reg__lane16_data   ) ,

    .reg__scntl__lane17_ready   ( reg__scntl__lane17_ready  ) ,
    .scntl__reg__lane17_valid   ( scntl__reg__lane17_valid  ) ,
    .scntl__reg__lane17_cntl    ( scntl__reg__lane17_cntl   ) ,
    .scntl__reg__lane17_data    ( scntl__reg__lane17_data   ) ,

    .reg__scntl__lane18_ready   ( reg__scntl__lane18_ready  ) ,
    .scntl__reg__lane18_valid   ( scntl__reg__lane18_valid  ) ,
    .scntl__reg__lane18_cntl    ( scntl__reg__lane18_cntl   ) ,
    .scntl__reg__lane18_data    ( scntl__reg__lane18_data   ) ,

    .reg__scntl__lane19_ready   ( reg__scntl__lane19_ready  ) ,
    .scntl__reg__lane19_valid   ( scntl__reg__lane19_valid  ) ,
    .scntl__reg__lane19_cntl    ( scntl__reg__lane19_cntl   ) ,
    .scntl__reg__lane19_data    ( scntl__reg__lane19_data   ) ,

    .reg__scntl__lane20_ready   ( reg__scntl__lane20_ready  ) ,
    .scntl__reg__lane20_valid   ( scntl__reg__lane20_valid  ) ,
    .scntl__reg__lane20_cntl    ( scntl__reg__lane20_cntl   ) ,
    .scntl__reg__lane20_data    ( scntl__reg__lane20_data   ) ,

    .reg__scntl__lane21_ready   ( reg__scntl__lane21_ready  ) ,
    .scntl__reg__lane21_valid   ( scntl__reg__lane21_valid  ) ,
    .scntl__reg__lane21_cntl    ( scntl__reg__lane21_cntl   ) ,
    .scntl__reg__lane21_data    ( scntl__reg__lane21_data   ) ,

    .reg__scntl__lane22_ready   ( reg__scntl__lane22_ready  ) ,
    .scntl__reg__lane22_valid   ( scntl__reg__lane22_valid  ) ,
    .scntl__reg__lane22_cntl    ( scntl__reg__lane22_cntl   ) ,
    .scntl__reg__lane22_data    ( scntl__reg__lane22_data   ) ,

    .reg__scntl__lane23_ready   ( reg__scntl__lane23_ready  ) ,
    .scntl__reg__lane23_valid   ( scntl__reg__lane23_valid  ) ,
    .scntl__reg__lane23_cntl    ( scntl__reg__lane23_cntl   ) ,
    .scntl__reg__lane23_data    ( scntl__reg__lane23_data   ) ,

    .reg__scntl__lane24_ready   ( reg__scntl__lane24_ready  ) ,
    .scntl__reg__lane24_valid   ( scntl__reg__lane24_valid  ) ,
    .scntl__reg__lane24_cntl    ( scntl__reg__lane24_cntl   ) ,
    .scntl__reg__lane24_data    ( scntl__reg__lane24_data   ) ,

    .reg__scntl__lane25_ready   ( reg__scntl__lane25_ready  ) ,
    .scntl__reg__lane25_valid   ( scntl__reg__lane25_valid  ) ,
    .scntl__reg__lane25_cntl    ( scntl__reg__lane25_cntl   ) ,
    .scntl__reg__lane25_data    ( scntl__reg__lane25_data   ) ,

    .reg__scntl__lane26_ready   ( reg__scntl__lane26_ready  ) ,
    .scntl__reg__lane26_valid   ( scntl__reg__lane26_valid  ) ,
    .scntl__reg__lane26_cntl    ( scntl__reg__lane26_cntl   ) ,
    .scntl__reg__lane26_data    ( scntl__reg__lane26_data   ) ,

    .reg__scntl__lane27_ready   ( reg__scntl__lane27_ready  ) ,
    .scntl__reg__lane27_valid   ( scntl__reg__lane27_valid  ) ,
    .scntl__reg__lane27_cntl    ( scntl__reg__lane27_cntl   ) ,
    .scntl__reg__lane27_data    ( scntl__reg__lane27_data   ) ,

    .reg__scntl__lane28_ready   ( reg__scntl__lane28_ready  ) ,
    .scntl__reg__lane28_valid   ( scntl__reg__lane28_valid  ) ,
    .scntl__reg__lane28_cntl    ( scntl__reg__lane28_cntl   ) ,
    .scntl__reg__lane28_data    ( scntl__reg__lane28_data   ) ,

    .reg__scntl__lane29_ready   ( reg__scntl__lane29_ready  ) ,
    .scntl__reg__lane29_valid   ( scntl__reg__lane29_valid  ) ,
    .scntl__reg__lane29_cntl    ( scntl__reg__lane29_cntl   ) ,
    .scntl__reg__lane29_data    ( scntl__reg__lane29_data   ) ,

    .reg__scntl__lane30_ready   ( reg__scntl__lane30_ready  ) ,
    .scntl__reg__lane30_valid   ( scntl__reg__lane30_valid  ) ,
    .scntl__reg__lane30_cntl    ( scntl__reg__lane30_cntl   ) ,
    .scntl__reg__lane30_data    ( scntl__reg__lane30_data   ) ,

    .reg__scntl__lane31_ready   ( reg__scntl__lane31_ready  ) ,
    .scntl__reg__lane31_valid   ( scntl__reg__lane31_valid  ) ,
    .scntl__reg__lane31_cntl    ( scntl__reg__lane31_cntl   ) ,
    .scntl__reg__lane31_data    ( scntl__reg__lane31_data   ) ,

