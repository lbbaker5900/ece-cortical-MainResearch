
    wire                                           stu__mgr0__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr0__cntl           ;
    wire                                           mgr0__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr0__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr0__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr0__oob_data       ;

    wire                                           stu__mgr1__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr1__cntl           ;
    wire                                           mgr1__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr1__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr1__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr1__oob_data       ;

    wire                                           stu__mgr2__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr2__cntl           ;
    wire                                           mgr2__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr2__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr2__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr2__oob_data       ;

    wire                                           stu__mgr3__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr3__cntl           ;
    wire                                           mgr3__stu__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr3__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr3__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr3__oob_data       ;

