
            fork                                                                                                                                  
                sys_operation_lane[0] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[0].Id[1]  =  0      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,0}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[0].put(sys_operation_lane[0])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[0];                                                                                                              
            join_none                                                                                                                             
            fork                                                                                                                                  
                sys_operation_lane[1] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[1].Id[1]  =  1      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,1}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[1].put(sys_operation_lane[1])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[1];                                                                                                              
            join_none                                                                                                                             
            fork                                                                                                                                  
                sys_operation_lane[2] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[2].Id[1]  =  2      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,2}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[2].put(sys_operation_lane[2])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[2];                                                                                                              
            join_none                                                                                                                             
            fork                                                                                                                                  
                sys_operation_lane[3] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[3].Id[1]  =  3      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,3}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[3].put(sys_operation_lane[3])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[3];                                                                                                              
            join_none                                                                                                                             
            fork                                                                                                                                  
                sys_operation_lane[4] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[4].Id[1]  =  4      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,4}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[4].put(sys_operation_lane[4])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[4];                                                                                                              
            join_none                                                                                                                             
            fork                                                                                                                                  
                sys_operation_lane[5] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[5].Id[1]  =  5      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,5}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[5].put(sys_operation_lane[5])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[5];                                                                                                              
            join_none                                                                                                                             
            fork                                                                                                                                  
                sys_operation_lane[6] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[6].Id[1]  =  6      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,6}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[6].put(sys_operation_lane[6])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[6];                                                                                                              
            join_none                                                                                                                             
            fork                                                                                                                                  
                sys_operation_lane[7] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[7].Id[1]  =  7      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,7}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[7].put(sys_operation_lane[7])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[7];                                                                                                              
            join_none                                                                                                                             
            fork                                                                                                                                  
                sys_operation_lane[8] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[8].Id[1]  =  8      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,8}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[8].put(sys_operation_lane[8])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[8];                                                                                                              
            join_none                                                                                                                             
            fork                                                                                                                                  
                sys_operation_lane[9] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[9].Id[1]  =  9      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,9}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[9].put(sys_operation_lane[9])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[9];                                                                                                              
            join_none                                                                                                                             
            fork                                                                                                                                  
                sys_operation_lane[10] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[10].Id[1]  =  10      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,10}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[10].put(sys_operation_lane[10])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[10];                                                                                                              
            join_none                                                                                                                             
            fork                                                                                                                                  
                sys_operation_lane[11] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[11].Id[1]  =  11      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,11}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[11].put(sys_operation_lane[11])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[11];                                                                                                              
            join_none                                                                                                                             
            fork                                                                                                                                  
                sys_operation_lane[12] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[12].Id[1]  =  12      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,12}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[12].put(sys_operation_lane[12])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[12];                                                                                                              
            join_none                                                                                                                             
            fork                                                                                                                                  
                sys_operation_lane[13] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[13].Id[1]  =  13      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,13}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[13].put(sys_operation_lane[13])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[13];                                                                                                              
            join_none                                                                                                                             
            fork                                                                                                                                  
                sys_operation_lane[14] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[14].Id[1]  =  14      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,14}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[14].put(sys_operation_lane[14])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[14];                                                                                                              
            join_none                                                                                                                             
            fork                                                                                                                                  
                sys_operation_lane[15] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[15].Id[1]  =  15      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,15}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[15].put(sys_operation_lane[15])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[15];                                                                                                              
            join_none                                                                                                                             
            fork                                                                                                                                  
                sys_operation_lane[16] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[16].Id[1]  =  16      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,16}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[16].put(sys_operation_lane[16])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[16];                                                                                                              
            join_none                                                                                                                             
            fork                                                                                                                                  
                sys_operation_lane[17] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[17].Id[1]  =  17      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,17}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[17].put(sys_operation_lane[17])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[17];                                                                                                              
            join_none                                                                                                                             
            fork                                                                                                                                  
                sys_operation_lane[18] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[18].Id[1]  =  18      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,18}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[18].put(sys_operation_lane[18])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[18];                                                                                                              
            join_none                                                                                                                             
            fork                                                                                                                                  
                sys_operation_lane[19] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[19].Id[1]  =  19      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,19}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[19].put(sys_operation_lane[19])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[19];                                                                                                              
            join_none                                                                                                                             
            fork                                                                                                                                  
                sys_operation_lane[20] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[20].Id[1]  =  20      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,20}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[20].put(sys_operation_lane[20])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[20];                                                                                                              
            join_none                                                                                                                             
            fork                                                                                                                                  
                sys_operation_lane[21] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[21].Id[1]  =  21      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,21}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[21].put(sys_operation_lane[21])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[21];                                                                                                              
            join_none                                                                                                                             
            fork                                                                                                                                  
                sys_operation_lane[22] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[22].Id[1]  =  22      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,22}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[22].put(sys_operation_lane[22])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[22];                                                                                                              
            join_none                                                                                                                             
            fork                                                                                                                                  
                sys_operation_lane[23] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[23].Id[1]  =  23      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,23}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[23].put(sys_operation_lane[23])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[23];                                                                                                              
            join_none                                                                                                                             
            fork                                                                                                                                  
                sys_operation_lane[24] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[24].Id[1]  =  24      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,24}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[24].put(sys_operation_lane[24])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[24];                                                                                                              
            join_none                                                                                                                             
            fork                                                                                                                                  
                sys_operation_lane[25] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[25].Id[1]  =  25      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,25}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[25].put(sys_operation_lane[25])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[25];                                                                                                              
            join_none                                                                                                                             
            fork                                                                                                                                  
                sys_operation_lane[26] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[26].Id[1]  =  26      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,26}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[26].put(sys_operation_lane[26])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[26];                                                                                                              
            join_none                                                                                                                             
            fork                                                                                                                                  
                sys_operation_lane[27] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[27].Id[1]  =  27      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,27}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[27].put(sys_operation_lane[27])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[27];                                                                                                              
            join_none                                                                                                                             
            fork                                                                                                                                  
                sys_operation_lane[28] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[28].Id[1]  =  28      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,28}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[28].put(sys_operation_lane[28])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[28];                                                                                                              
            join_none                                                                                                                             
            fork                                                                                                                                  
                sys_operation_lane[29] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[29].Id[1]  =  29      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,29}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[29].put(sys_operation_lane[29])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[29];                                                                                                              
            join_none                                                                                                                             
            fork                                                                                                                                  
                sys_operation_lane[30] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[30].Id[1]  =  30      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,30}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[30].put(sys_operation_lane[30])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[30];                                                                                                              
            join_none                                                                                                                             
            fork                                                                                                                                  
                sys_operation_lane[31] = sys_operation_mgr.copy() ; // deep copy creates new operand arrays                                      
                sys_operation_lane[31].Id[1]  =  31      ;  // set lane for address generation                                                  
                                                                                                                                                  
                // Send to driver                                                                                                                 
                //$display("@%0t:%s:%0d:LEE: sys_operation_mgr : {%0d,31}:%h\n", $time, `__FILE__, `__LINE__, Id, sys_operation_mgr);            
                mgr2gen[31].put(sys_operation_lane[31])                    ;                                                                    
                                                                                                                                                  
                // now wait for generator                                                                                                         
                //sys_operation.displayOperation();                                                                                               
                @mgr2gen_ack[31];                                                                                                              
            join_none                                                                                                                             
