
  // Common (Scalar) Register(s)                
  assign   simd__cntl__rs0  = cntl__simd__rs0 ;
  assign   simd__cntl__rs1  = cntl__simd__rs1 ;

  // Lane Register(s)                
// Lane 0                 
  assign  simd__cntl__lane_r128  [0]   =   cntl__simd__lane_r128  [0]  ;
  assign  simd__cntl__lane_r129  [0]   =   cntl__simd__lane_r129  [0]  ;
  assign  simd__cntl__lane_r130  [0]   =   cntl__simd__lane_r130  [0]  ;
  assign  simd__cntl__lane_r131  [0]   =   cntl__simd__lane_r131  [0]  ;
  assign  simd__cntl__lane_r132  [0]   =   cntl__simd__lane_r132  [0]  ;
  assign  simd__cntl__lane_r133  [0]   =   cntl__simd__lane_r133  [0]  ;
  assign  simd__cntl__lane_r134  [0]   =   cntl__simd__lane_r134  [0]  ;
  assign  simd__cntl__lane_r135  [0]   =   cntl__simd__lane_r135  [0]  ;

// Lane 1                 
  assign  simd__cntl__lane_r128  [1]   =   cntl__simd__lane_r128  [1]  ;
  assign  simd__cntl__lane_r129  [1]   =   cntl__simd__lane_r129  [1]  ;
  assign  simd__cntl__lane_r130  [1]   =   cntl__simd__lane_r130  [1]  ;
  assign  simd__cntl__lane_r131  [1]   =   cntl__simd__lane_r131  [1]  ;
  assign  simd__cntl__lane_r132  [1]   =   cntl__simd__lane_r132  [1]  ;
  assign  simd__cntl__lane_r133  [1]   =   cntl__simd__lane_r133  [1]  ;
  assign  simd__cntl__lane_r134  [1]   =   cntl__simd__lane_r134  [1]  ;
  assign  simd__cntl__lane_r135  [1]   =   cntl__simd__lane_r135  [1]  ;

// Lane 2                 
  assign  simd__cntl__lane_r128  [2]   =   cntl__simd__lane_r128  [2]  ;
  assign  simd__cntl__lane_r129  [2]   =   cntl__simd__lane_r129  [2]  ;
  assign  simd__cntl__lane_r130  [2]   =   cntl__simd__lane_r130  [2]  ;
  assign  simd__cntl__lane_r131  [2]   =   cntl__simd__lane_r131  [2]  ;
  assign  simd__cntl__lane_r132  [2]   =   cntl__simd__lane_r132  [2]  ;
  assign  simd__cntl__lane_r133  [2]   =   cntl__simd__lane_r133  [2]  ;
  assign  simd__cntl__lane_r134  [2]   =   cntl__simd__lane_r134  [2]  ;
  assign  simd__cntl__lane_r135  [2]   =   cntl__simd__lane_r135  [2]  ;

// Lane 3                 
  assign  simd__cntl__lane_r128  [3]   =   cntl__simd__lane_r128  [3]  ;
  assign  simd__cntl__lane_r129  [3]   =   cntl__simd__lane_r129  [3]  ;
  assign  simd__cntl__lane_r130  [3]   =   cntl__simd__lane_r130  [3]  ;
  assign  simd__cntl__lane_r131  [3]   =   cntl__simd__lane_r131  [3]  ;
  assign  simd__cntl__lane_r132  [3]   =   cntl__simd__lane_r132  [3]  ;
  assign  simd__cntl__lane_r133  [3]   =   cntl__simd__lane_r133  [3]  ;
  assign  simd__cntl__lane_r134  [3]   =   cntl__simd__lane_r134  [3]  ;
  assign  simd__cntl__lane_r135  [3]   =   cntl__simd__lane_r135  [3]  ;

// Lane 4                 
  assign  simd__cntl__lane_r128  [4]   =   cntl__simd__lane_r128  [4]  ;
  assign  simd__cntl__lane_r129  [4]   =   cntl__simd__lane_r129  [4]  ;
  assign  simd__cntl__lane_r130  [4]   =   cntl__simd__lane_r130  [4]  ;
  assign  simd__cntl__lane_r131  [4]   =   cntl__simd__lane_r131  [4]  ;
  assign  simd__cntl__lane_r132  [4]   =   cntl__simd__lane_r132  [4]  ;
  assign  simd__cntl__lane_r133  [4]   =   cntl__simd__lane_r133  [4]  ;
  assign  simd__cntl__lane_r134  [4]   =   cntl__simd__lane_r134  [4]  ;
  assign  simd__cntl__lane_r135  [4]   =   cntl__simd__lane_r135  [4]  ;

// Lane 5                 
  assign  simd__cntl__lane_r128  [5]   =   cntl__simd__lane_r128  [5]  ;
  assign  simd__cntl__lane_r129  [5]   =   cntl__simd__lane_r129  [5]  ;
  assign  simd__cntl__lane_r130  [5]   =   cntl__simd__lane_r130  [5]  ;
  assign  simd__cntl__lane_r131  [5]   =   cntl__simd__lane_r131  [5]  ;
  assign  simd__cntl__lane_r132  [5]   =   cntl__simd__lane_r132  [5]  ;
  assign  simd__cntl__lane_r133  [5]   =   cntl__simd__lane_r133  [5]  ;
  assign  simd__cntl__lane_r134  [5]   =   cntl__simd__lane_r134  [5]  ;
  assign  simd__cntl__lane_r135  [5]   =   cntl__simd__lane_r135  [5]  ;

// Lane 6                 
  assign  simd__cntl__lane_r128  [6]   =   cntl__simd__lane_r128  [6]  ;
  assign  simd__cntl__lane_r129  [6]   =   cntl__simd__lane_r129  [6]  ;
  assign  simd__cntl__lane_r130  [6]   =   cntl__simd__lane_r130  [6]  ;
  assign  simd__cntl__lane_r131  [6]   =   cntl__simd__lane_r131  [6]  ;
  assign  simd__cntl__lane_r132  [6]   =   cntl__simd__lane_r132  [6]  ;
  assign  simd__cntl__lane_r133  [6]   =   cntl__simd__lane_r133  [6]  ;
  assign  simd__cntl__lane_r134  [6]   =   cntl__simd__lane_r134  [6]  ;
  assign  simd__cntl__lane_r135  [6]   =   cntl__simd__lane_r135  [6]  ;

// Lane 7                 
  assign  simd__cntl__lane_r128  [7]   =   cntl__simd__lane_r128  [7]  ;
  assign  simd__cntl__lane_r129  [7]   =   cntl__simd__lane_r129  [7]  ;
  assign  simd__cntl__lane_r130  [7]   =   cntl__simd__lane_r130  [7]  ;
  assign  simd__cntl__lane_r131  [7]   =   cntl__simd__lane_r131  [7]  ;
  assign  simd__cntl__lane_r132  [7]   =   cntl__simd__lane_r132  [7]  ;
  assign  simd__cntl__lane_r133  [7]   =   cntl__simd__lane_r133  [7]  ;
  assign  simd__cntl__lane_r134  [7]   =   cntl__simd__lane_r134  [7]  ;
  assign  simd__cntl__lane_r135  [7]   =   cntl__simd__lane_r135  [7]  ;

// Lane 8                 
  assign  simd__cntl__lane_r128  [8]   =   cntl__simd__lane_r128  [8]  ;
  assign  simd__cntl__lane_r129  [8]   =   cntl__simd__lane_r129  [8]  ;
  assign  simd__cntl__lane_r130  [8]   =   cntl__simd__lane_r130  [8]  ;
  assign  simd__cntl__lane_r131  [8]   =   cntl__simd__lane_r131  [8]  ;
  assign  simd__cntl__lane_r132  [8]   =   cntl__simd__lane_r132  [8]  ;
  assign  simd__cntl__lane_r133  [8]   =   cntl__simd__lane_r133  [8]  ;
  assign  simd__cntl__lane_r134  [8]   =   cntl__simd__lane_r134  [8]  ;
  assign  simd__cntl__lane_r135  [8]   =   cntl__simd__lane_r135  [8]  ;

// Lane 9                 
  assign  simd__cntl__lane_r128  [9]   =   cntl__simd__lane_r128  [9]  ;
  assign  simd__cntl__lane_r129  [9]   =   cntl__simd__lane_r129  [9]  ;
  assign  simd__cntl__lane_r130  [9]   =   cntl__simd__lane_r130  [9]  ;
  assign  simd__cntl__lane_r131  [9]   =   cntl__simd__lane_r131  [9]  ;
  assign  simd__cntl__lane_r132  [9]   =   cntl__simd__lane_r132  [9]  ;
  assign  simd__cntl__lane_r133  [9]   =   cntl__simd__lane_r133  [9]  ;
  assign  simd__cntl__lane_r134  [9]   =   cntl__simd__lane_r134  [9]  ;
  assign  simd__cntl__lane_r135  [9]   =   cntl__simd__lane_r135  [9]  ;

// Lane 10                 
  assign  simd__cntl__lane_r128  [10]   =   cntl__simd__lane_r128  [10]  ;
  assign  simd__cntl__lane_r129  [10]   =   cntl__simd__lane_r129  [10]  ;
  assign  simd__cntl__lane_r130  [10]   =   cntl__simd__lane_r130  [10]  ;
  assign  simd__cntl__lane_r131  [10]   =   cntl__simd__lane_r131  [10]  ;
  assign  simd__cntl__lane_r132  [10]   =   cntl__simd__lane_r132  [10]  ;
  assign  simd__cntl__lane_r133  [10]   =   cntl__simd__lane_r133  [10]  ;
  assign  simd__cntl__lane_r134  [10]   =   cntl__simd__lane_r134  [10]  ;
  assign  simd__cntl__lane_r135  [10]   =   cntl__simd__lane_r135  [10]  ;

// Lane 11                 
  assign  simd__cntl__lane_r128  [11]   =   cntl__simd__lane_r128  [11]  ;
  assign  simd__cntl__lane_r129  [11]   =   cntl__simd__lane_r129  [11]  ;
  assign  simd__cntl__lane_r130  [11]   =   cntl__simd__lane_r130  [11]  ;
  assign  simd__cntl__lane_r131  [11]   =   cntl__simd__lane_r131  [11]  ;
  assign  simd__cntl__lane_r132  [11]   =   cntl__simd__lane_r132  [11]  ;
  assign  simd__cntl__lane_r133  [11]   =   cntl__simd__lane_r133  [11]  ;
  assign  simd__cntl__lane_r134  [11]   =   cntl__simd__lane_r134  [11]  ;
  assign  simd__cntl__lane_r135  [11]   =   cntl__simd__lane_r135  [11]  ;

// Lane 12                 
  assign  simd__cntl__lane_r128  [12]   =   cntl__simd__lane_r128  [12]  ;
  assign  simd__cntl__lane_r129  [12]   =   cntl__simd__lane_r129  [12]  ;
  assign  simd__cntl__lane_r130  [12]   =   cntl__simd__lane_r130  [12]  ;
  assign  simd__cntl__lane_r131  [12]   =   cntl__simd__lane_r131  [12]  ;
  assign  simd__cntl__lane_r132  [12]   =   cntl__simd__lane_r132  [12]  ;
  assign  simd__cntl__lane_r133  [12]   =   cntl__simd__lane_r133  [12]  ;
  assign  simd__cntl__lane_r134  [12]   =   cntl__simd__lane_r134  [12]  ;
  assign  simd__cntl__lane_r135  [12]   =   cntl__simd__lane_r135  [12]  ;

// Lane 13                 
  assign  simd__cntl__lane_r128  [13]   =   cntl__simd__lane_r128  [13]  ;
  assign  simd__cntl__lane_r129  [13]   =   cntl__simd__lane_r129  [13]  ;
  assign  simd__cntl__lane_r130  [13]   =   cntl__simd__lane_r130  [13]  ;
  assign  simd__cntl__lane_r131  [13]   =   cntl__simd__lane_r131  [13]  ;
  assign  simd__cntl__lane_r132  [13]   =   cntl__simd__lane_r132  [13]  ;
  assign  simd__cntl__lane_r133  [13]   =   cntl__simd__lane_r133  [13]  ;
  assign  simd__cntl__lane_r134  [13]   =   cntl__simd__lane_r134  [13]  ;
  assign  simd__cntl__lane_r135  [13]   =   cntl__simd__lane_r135  [13]  ;

// Lane 14                 
  assign  simd__cntl__lane_r128  [14]   =   cntl__simd__lane_r128  [14]  ;
  assign  simd__cntl__lane_r129  [14]   =   cntl__simd__lane_r129  [14]  ;
  assign  simd__cntl__lane_r130  [14]   =   cntl__simd__lane_r130  [14]  ;
  assign  simd__cntl__lane_r131  [14]   =   cntl__simd__lane_r131  [14]  ;
  assign  simd__cntl__lane_r132  [14]   =   cntl__simd__lane_r132  [14]  ;
  assign  simd__cntl__lane_r133  [14]   =   cntl__simd__lane_r133  [14]  ;
  assign  simd__cntl__lane_r134  [14]   =   cntl__simd__lane_r134  [14]  ;
  assign  simd__cntl__lane_r135  [14]   =   cntl__simd__lane_r135  [14]  ;

// Lane 15                 
  assign  simd__cntl__lane_r128  [15]   =   cntl__simd__lane_r128  [15]  ;
  assign  simd__cntl__lane_r129  [15]   =   cntl__simd__lane_r129  [15]  ;
  assign  simd__cntl__lane_r130  [15]   =   cntl__simd__lane_r130  [15]  ;
  assign  simd__cntl__lane_r131  [15]   =   cntl__simd__lane_r131  [15]  ;
  assign  simd__cntl__lane_r132  [15]   =   cntl__simd__lane_r132  [15]  ;
  assign  simd__cntl__lane_r133  [15]   =   cntl__simd__lane_r133  [15]  ;
  assign  simd__cntl__lane_r134  [15]   =   cntl__simd__lane_r134  [15]  ;
  assign  simd__cntl__lane_r135  [15]   =   cntl__simd__lane_r135  [15]  ;

// Lane 16                 
  assign  simd__cntl__lane_r128  [16]   =   cntl__simd__lane_r128  [16]  ;
  assign  simd__cntl__lane_r129  [16]   =   cntl__simd__lane_r129  [16]  ;
  assign  simd__cntl__lane_r130  [16]   =   cntl__simd__lane_r130  [16]  ;
  assign  simd__cntl__lane_r131  [16]   =   cntl__simd__lane_r131  [16]  ;
  assign  simd__cntl__lane_r132  [16]   =   cntl__simd__lane_r132  [16]  ;
  assign  simd__cntl__lane_r133  [16]   =   cntl__simd__lane_r133  [16]  ;
  assign  simd__cntl__lane_r134  [16]   =   cntl__simd__lane_r134  [16]  ;
  assign  simd__cntl__lane_r135  [16]   =   cntl__simd__lane_r135  [16]  ;

// Lane 17                 
  assign  simd__cntl__lane_r128  [17]   =   cntl__simd__lane_r128  [17]  ;
  assign  simd__cntl__lane_r129  [17]   =   cntl__simd__lane_r129  [17]  ;
  assign  simd__cntl__lane_r130  [17]   =   cntl__simd__lane_r130  [17]  ;
  assign  simd__cntl__lane_r131  [17]   =   cntl__simd__lane_r131  [17]  ;
  assign  simd__cntl__lane_r132  [17]   =   cntl__simd__lane_r132  [17]  ;
  assign  simd__cntl__lane_r133  [17]   =   cntl__simd__lane_r133  [17]  ;
  assign  simd__cntl__lane_r134  [17]   =   cntl__simd__lane_r134  [17]  ;
  assign  simd__cntl__lane_r135  [17]   =   cntl__simd__lane_r135  [17]  ;

// Lane 18                 
  assign  simd__cntl__lane_r128  [18]   =   cntl__simd__lane_r128  [18]  ;
  assign  simd__cntl__lane_r129  [18]   =   cntl__simd__lane_r129  [18]  ;
  assign  simd__cntl__lane_r130  [18]   =   cntl__simd__lane_r130  [18]  ;
  assign  simd__cntl__lane_r131  [18]   =   cntl__simd__lane_r131  [18]  ;
  assign  simd__cntl__lane_r132  [18]   =   cntl__simd__lane_r132  [18]  ;
  assign  simd__cntl__lane_r133  [18]   =   cntl__simd__lane_r133  [18]  ;
  assign  simd__cntl__lane_r134  [18]   =   cntl__simd__lane_r134  [18]  ;
  assign  simd__cntl__lane_r135  [18]   =   cntl__simd__lane_r135  [18]  ;

// Lane 19                 
  assign  simd__cntl__lane_r128  [19]   =   cntl__simd__lane_r128  [19]  ;
  assign  simd__cntl__lane_r129  [19]   =   cntl__simd__lane_r129  [19]  ;
  assign  simd__cntl__lane_r130  [19]   =   cntl__simd__lane_r130  [19]  ;
  assign  simd__cntl__lane_r131  [19]   =   cntl__simd__lane_r131  [19]  ;
  assign  simd__cntl__lane_r132  [19]   =   cntl__simd__lane_r132  [19]  ;
  assign  simd__cntl__lane_r133  [19]   =   cntl__simd__lane_r133  [19]  ;
  assign  simd__cntl__lane_r134  [19]   =   cntl__simd__lane_r134  [19]  ;
  assign  simd__cntl__lane_r135  [19]   =   cntl__simd__lane_r135  [19]  ;

// Lane 20                 
  assign  simd__cntl__lane_r128  [20]   =   cntl__simd__lane_r128  [20]  ;
  assign  simd__cntl__lane_r129  [20]   =   cntl__simd__lane_r129  [20]  ;
  assign  simd__cntl__lane_r130  [20]   =   cntl__simd__lane_r130  [20]  ;
  assign  simd__cntl__lane_r131  [20]   =   cntl__simd__lane_r131  [20]  ;
  assign  simd__cntl__lane_r132  [20]   =   cntl__simd__lane_r132  [20]  ;
  assign  simd__cntl__lane_r133  [20]   =   cntl__simd__lane_r133  [20]  ;
  assign  simd__cntl__lane_r134  [20]   =   cntl__simd__lane_r134  [20]  ;
  assign  simd__cntl__lane_r135  [20]   =   cntl__simd__lane_r135  [20]  ;

// Lane 21                 
  assign  simd__cntl__lane_r128  [21]   =   cntl__simd__lane_r128  [21]  ;
  assign  simd__cntl__lane_r129  [21]   =   cntl__simd__lane_r129  [21]  ;
  assign  simd__cntl__lane_r130  [21]   =   cntl__simd__lane_r130  [21]  ;
  assign  simd__cntl__lane_r131  [21]   =   cntl__simd__lane_r131  [21]  ;
  assign  simd__cntl__lane_r132  [21]   =   cntl__simd__lane_r132  [21]  ;
  assign  simd__cntl__lane_r133  [21]   =   cntl__simd__lane_r133  [21]  ;
  assign  simd__cntl__lane_r134  [21]   =   cntl__simd__lane_r134  [21]  ;
  assign  simd__cntl__lane_r135  [21]   =   cntl__simd__lane_r135  [21]  ;

// Lane 22                 
  assign  simd__cntl__lane_r128  [22]   =   cntl__simd__lane_r128  [22]  ;
  assign  simd__cntl__lane_r129  [22]   =   cntl__simd__lane_r129  [22]  ;
  assign  simd__cntl__lane_r130  [22]   =   cntl__simd__lane_r130  [22]  ;
  assign  simd__cntl__lane_r131  [22]   =   cntl__simd__lane_r131  [22]  ;
  assign  simd__cntl__lane_r132  [22]   =   cntl__simd__lane_r132  [22]  ;
  assign  simd__cntl__lane_r133  [22]   =   cntl__simd__lane_r133  [22]  ;
  assign  simd__cntl__lane_r134  [22]   =   cntl__simd__lane_r134  [22]  ;
  assign  simd__cntl__lane_r135  [22]   =   cntl__simd__lane_r135  [22]  ;

// Lane 23                 
  assign  simd__cntl__lane_r128  [23]   =   cntl__simd__lane_r128  [23]  ;
  assign  simd__cntl__lane_r129  [23]   =   cntl__simd__lane_r129  [23]  ;
  assign  simd__cntl__lane_r130  [23]   =   cntl__simd__lane_r130  [23]  ;
  assign  simd__cntl__lane_r131  [23]   =   cntl__simd__lane_r131  [23]  ;
  assign  simd__cntl__lane_r132  [23]   =   cntl__simd__lane_r132  [23]  ;
  assign  simd__cntl__lane_r133  [23]   =   cntl__simd__lane_r133  [23]  ;
  assign  simd__cntl__lane_r134  [23]   =   cntl__simd__lane_r134  [23]  ;
  assign  simd__cntl__lane_r135  [23]   =   cntl__simd__lane_r135  [23]  ;

// Lane 24                 
  assign  simd__cntl__lane_r128  [24]   =   cntl__simd__lane_r128  [24]  ;
  assign  simd__cntl__lane_r129  [24]   =   cntl__simd__lane_r129  [24]  ;
  assign  simd__cntl__lane_r130  [24]   =   cntl__simd__lane_r130  [24]  ;
  assign  simd__cntl__lane_r131  [24]   =   cntl__simd__lane_r131  [24]  ;
  assign  simd__cntl__lane_r132  [24]   =   cntl__simd__lane_r132  [24]  ;
  assign  simd__cntl__lane_r133  [24]   =   cntl__simd__lane_r133  [24]  ;
  assign  simd__cntl__lane_r134  [24]   =   cntl__simd__lane_r134  [24]  ;
  assign  simd__cntl__lane_r135  [24]   =   cntl__simd__lane_r135  [24]  ;

// Lane 25                 
  assign  simd__cntl__lane_r128  [25]   =   cntl__simd__lane_r128  [25]  ;
  assign  simd__cntl__lane_r129  [25]   =   cntl__simd__lane_r129  [25]  ;
  assign  simd__cntl__lane_r130  [25]   =   cntl__simd__lane_r130  [25]  ;
  assign  simd__cntl__lane_r131  [25]   =   cntl__simd__lane_r131  [25]  ;
  assign  simd__cntl__lane_r132  [25]   =   cntl__simd__lane_r132  [25]  ;
  assign  simd__cntl__lane_r133  [25]   =   cntl__simd__lane_r133  [25]  ;
  assign  simd__cntl__lane_r134  [25]   =   cntl__simd__lane_r134  [25]  ;
  assign  simd__cntl__lane_r135  [25]   =   cntl__simd__lane_r135  [25]  ;

// Lane 26                 
  assign  simd__cntl__lane_r128  [26]   =   cntl__simd__lane_r128  [26]  ;
  assign  simd__cntl__lane_r129  [26]   =   cntl__simd__lane_r129  [26]  ;
  assign  simd__cntl__lane_r130  [26]   =   cntl__simd__lane_r130  [26]  ;
  assign  simd__cntl__lane_r131  [26]   =   cntl__simd__lane_r131  [26]  ;
  assign  simd__cntl__lane_r132  [26]   =   cntl__simd__lane_r132  [26]  ;
  assign  simd__cntl__lane_r133  [26]   =   cntl__simd__lane_r133  [26]  ;
  assign  simd__cntl__lane_r134  [26]   =   cntl__simd__lane_r134  [26]  ;
  assign  simd__cntl__lane_r135  [26]   =   cntl__simd__lane_r135  [26]  ;

// Lane 27                 
  assign  simd__cntl__lane_r128  [27]   =   cntl__simd__lane_r128  [27]  ;
  assign  simd__cntl__lane_r129  [27]   =   cntl__simd__lane_r129  [27]  ;
  assign  simd__cntl__lane_r130  [27]   =   cntl__simd__lane_r130  [27]  ;
  assign  simd__cntl__lane_r131  [27]   =   cntl__simd__lane_r131  [27]  ;
  assign  simd__cntl__lane_r132  [27]   =   cntl__simd__lane_r132  [27]  ;
  assign  simd__cntl__lane_r133  [27]   =   cntl__simd__lane_r133  [27]  ;
  assign  simd__cntl__lane_r134  [27]   =   cntl__simd__lane_r134  [27]  ;
  assign  simd__cntl__lane_r135  [27]   =   cntl__simd__lane_r135  [27]  ;

// Lane 28                 
  assign  simd__cntl__lane_r128  [28]   =   cntl__simd__lane_r128  [28]  ;
  assign  simd__cntl__lane_r129  [28]   =   cntl__simd__lane_r129  [28]  ;
  assign  simd__cntl__lane_r130  [28]   =   cntl__simd__lane_r130  [28]  ;
  assign  simd__cntl__lane_r131  [28]   =   cntl__simd__lane_r131  [28]  ;
  assign  simd__cntl__lane_r132  [28]   =   cntl__simd__lane_r132  [28]  ;
  assign  simd__cntl__lane_r133  [28]   =   cntl__simd__lane_r133  [28]  ;
  assign  simd__cntl__lane_r134  [28]   =   cntl__simd__lane_r134  [28]  ;
  assign  simd__cntl__lane_r135  [28]   =   cntl__simd__lane_r135  [28]  ;

// Lane 29                 
  assign  simd__cntl__lane_r128  [29]   =   cntl__simd__lane_r128  [29]  ;
  assign  simd__cntl__lane_r129  [29]   =   cntl__simd__lane_r129  [29]  ;
  assign  simd__cntl__lane_r130  [29]   =   cntl__simd__lane_r130  [29]  ;
  assign  simd__cntl__lane_r131  [29]   =   cntl__simd__lane_r131  [29]  ;
  assign  simd__cntl__lane_r132  [29]   =   cntl__simd__lane_r132  [29]  ;
  assign  simd__cntl__lane_r133  [29]   =   cntl__simd__lane_r133  [29]  ;
  assign  simd__cntl__lane_r134  [29]   =   cntl__simd__lane_r134  [29]  ;
  assign  simd__cntl__lane_r135  [29]   =   cntl__simd__lane_r135  [29]  ;

// Lane 30                 
  assign  simd__cntl__lane_r128  [30]   =   cntl__simd__lane_r128  [30]  ;
  assign  simd__cntl__lane_r129  [30]   =   cntl__simd__lane_r129  [30]  ;
  assign  simd__cntl__lane_r130  [30]   =   cntl__simd__lane_r130  [30]  ;
  assign  simd__cntl__lane_r131  [30]   =   cntl__simd__lane_r131  [30]  ;
  assign  simd__cntl__lane_r132  [30]   =   cntl__simd__lane_r132  [30]  ;
  assign  simd__cntl__lane_r133  [30]   =   cntl__simd__lane_r133  [30]  ;
  assign  simd__cntl__lane_r134  [30]   =   cntl__simd__lane_r134  [30]  ;
  assign  simd__cntl__lane_r135  [30]   =   cntl__simd__lane_r135  [30]  ;

// Lane 31                 
  assign  simd__cntl__lane_r128  [31]   =   cntl__simd__lane_r128  [31]  ;
  assign  simd__cntl__lane_r129  [31]   =   cntl__simd__lane_r129  [31]  ;
  assign  simd__cntl__lane_r130  [31]   =   cntl__simd__lane_r130  [31]  ;
  assign  simd__cntl__lane_r131  [31]   =   cntl__simd__lane_r131  [31]  ;
  assign  simd__cntl__lane_r132  [31]   =   cntl__simd__lane_r132  [31]  ;
  assign  simd__cntl__lane_r133  [31]   =   cntl__simd__lane_r133  [31]  ;
  assign  simd__cntl__lane_r134  [31]   =   cntl__simd__lane_r134  [31]  ;
  assign  simd__cntl__lane_r135  [31]   =   cntl__simd__lane_r135  [31]  ;

